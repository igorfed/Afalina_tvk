-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_mux 

-- ============================================================
-- File Name: MUX_REG.vhd
-- Megafunction Name(s):
-- 			lpm_mux
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 7.2 Build 151 09/26/2007 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2007 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY MUX_REG IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data100x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data101x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data102x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data103x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data104x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data105x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data106x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data107x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data108x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data109x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data10x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data110x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data111x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data112x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data113x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data114x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data115x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data116x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data117x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data118x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data119x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data11x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data120x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data121x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data122x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data123x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data124x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data125x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data126x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data127x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data128x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data129x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data12x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data130x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data131x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data132x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data133x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data134x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data135x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data136x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data137x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data138x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data139x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data13x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data140x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data141x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data142x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data143x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data144x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data145x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data146x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data147x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data148x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data149x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data14x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data150x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data151x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data152x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data153x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data154x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data155x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data156x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data157x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data158x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data159x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data15x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data160x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data161x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data162x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data163x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data164x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data165x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data166x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data167x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data168x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data169x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data16x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data170x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data171x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data172x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data173x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data174x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data175x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data176x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data177x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data178x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data179x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data17x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data180x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data181x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data182x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data183x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data184x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data185x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data186x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data187x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data188x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data189x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data18x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data190x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data191x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data192x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data193x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data194x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data195x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data196x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data197x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data198x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data199x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data19x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data200x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data201x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data202x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data203x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data204x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data205x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data206x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data207x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data208x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data209x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data20x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data210x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data211x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data212x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data213x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data214x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data215x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data216x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data217x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data218x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data219x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data21x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data220x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data221x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data222x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data223x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data224x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data225x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data226x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data227x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data228x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data229x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data22x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data230x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data231x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data232x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data233x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data234x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data235x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data236x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data237x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data238x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data239x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data23x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data240x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data241x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data242x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data243x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data244x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data245x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data246x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data247x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data248x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data249x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data24x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data250x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data251x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data252x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data253x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data254x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data255x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data25x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data26x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data27x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data28x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data29x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data30x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data31x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data32x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data33x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data34x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data35x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data36x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data37x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data38x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data39x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data40x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data41x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data42x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data43x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data44x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data45x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data46x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data47x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data48x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data49x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data50x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data51x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data52x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data53x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data54x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data55x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data56x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data57x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data58x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data59x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data60x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data61x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data62x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data63x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data64x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data65x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data66x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data67x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data68x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data69x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data70x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data71x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data72x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data73x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data74x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data75x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data76x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data77x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data78x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data79x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data80x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data81x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data82x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data83x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data84x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data85x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data86x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data87x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data88x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data89x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data8x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data90x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data91x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data92x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data93x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data94x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data95x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data96x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data97x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data98x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data99x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		data9x		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END MUX_REG;


ARCHITECTURE SYN OF mux_reg IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_2D (255 DOWNTO 0, 7 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire18	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire19	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire20	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire21	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire22	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire23	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire24	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire25	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire26	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire27	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire28	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire29	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire30	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire31	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire32	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire33	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire34	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire35	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire36	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire37	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire38	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire39	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire40	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire41	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire42	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire43	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire44	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire45	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire46	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire47	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire48	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire49	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire50	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire51	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire52	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire53	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire54	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire55	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire56	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire57	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire58	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire59	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire60	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire61	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire62	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire63	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire64	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire65	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire66	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire67	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire68	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire69	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire70	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire71	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire72	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire73	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire74	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire75	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire76	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire77	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire78	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire79	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire80	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire81	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire82	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire83	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire84	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire85	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire86	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire87	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire88	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire89	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire90	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire91	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire92	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire93	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire94	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire95	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire96	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire97	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire98	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire99	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire100	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire101	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire102	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire103	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire104	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire105	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire106	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire107	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire108	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire109	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire110	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire111	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire112	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire113	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire114	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire115	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire116	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire117	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire118	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire119	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire120	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire121	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire122	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire123	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire124	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire125	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire126	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire127	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire128	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire129	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire130	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire131	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire132	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire133	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire134	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire135	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire136	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire137	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire138	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire139	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire140	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire141	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire142	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire143	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire144	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire145	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire146	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire147	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire148	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire149	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire150	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire151	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire152	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire153	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire154	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire155	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire156	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire157	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire158	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire159	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire160	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire161	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire162	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire163	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire164	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire165	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire166	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire167	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire168	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire169	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire170	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire171	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire172	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire173	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire174	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire175	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire176	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire177	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire178	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire179	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire180	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire181	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire182	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire183	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire184	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire185	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire186	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire187	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire188	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire189	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire190	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire191	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire192	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire193	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire194	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire195	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire196	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire197	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire198	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire199	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire200	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire201	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire202	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire203	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire204	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire205	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire206	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire207	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire208	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire209	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire210	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire211	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire212	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire213	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire214	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire215	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire216	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire217	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire218	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire219	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire220	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire221	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire222	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire223	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire224	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire225	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire226	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire227	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire228	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire229	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire230	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire231	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire232	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire233	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire234	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire235	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire236	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire237	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire238	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire239	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire240	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire241	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire242	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire243	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire244	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire245	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire246	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire247	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire248	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire249	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire250	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire251	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire252	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire253	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire254	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire255	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire256	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire257	: STD_LOGIC_VECTOR (7 DOWNTO 0);

BEGIN
	sub_wire257    <= data0x(7 DOWNTO 0);
	sub_wire256    <= data1x(7 DOWNTO 0);
	sub_wire255    <= data2x(7 DOWNTO 0);
	sub_wire254    <= data3x(7 DOWNTO 0);
	sub_wire253    <= data4x(7 DOWNTO 0);
	sub_wire252    <= data5x(7 DOWNTO 0);
	sub_wire251    <= data6x(7 DOWNTO 0);
	sub_wire250    <= data7x(7 DOWNTO 0);
	sub_wire249    <= data8x(7 DOWNTO 0);
	sub_wire248    <= data9x(7 DOWNTO 0);
	sub_wire247    <= data10x(7 DOWNTO 0);
	sub_wire246    <= data11x(7 DOWNTO 0);
	sub_wire245    <= data12x(7 DOWNTO 0);
	sub_wire244    <= data13x(7 DOWNTO 0);
	sub_wire243    <= data14x(7 DOWNTO 0);
	sub_wire242    <= data15x(7 DOWNTO 0);
	sub_wire241    <= data16x(7 DOWNTO 0);
	sub_wire240    <= data17x(7 DOWNTO 0);
	sub_wire239    <= data18x(7 DOWNTO 0);
	sub_wire238    <= data19x(7 DOWNTO 0);
	sub_wire237    <= data20x(7 DOWNTO 0);
	sub_wire236    <= data21x(7 DOWNTO 0);
	sub_wire235    <= data22x(7 DOWNTO 0);
	sub_wire234    <= data23x(7 DOWNTO 0);
	sub_wire233    <= data24x(7 DOWNTO 0);
	sub_wire232    <= data25x(7 DOWNTO 0);
	sub_wire231    <= data26x(7 DOWNTO 0);
	sub_wire230    <= data27x(7 DOWNTO 0);
	sub_wire229    <= data28x(7 DOWNTO 0);
	sub_wire228    <= data29x(7 DOWNTO 0);
	sub_wire227    <= data30x(7 DOWNTO 0);
	sub_wire226    <= data31x(7 DOWNTO 0);
	sub_wire225    <= data32x(7 DOWNTO 0);
	sub_wire224    <= data33x(7 DOWNTO 0);
	sub_wire223    <= data34x(7 DOWNTO 0);
	sub_wire222    <= data35x(7 DOWNTO 0);
	sub_wire221    <= data36x(7 DOWNTO 0);
	sub_wire220    <= data37x(7 DOWNTO 0);
	sub_wire219    <= data38x(7 DOWNTO 0);
	sub_wire218    <= data39x(7 DOWNTO 0);
	sub_wire217    <= data40x(7 DOWNTO 0);
	sub_wire216    <= data41x(7 DOWNTO 0);
	sub_wire215    <= data42x(7 DOWNTO 0);
	sub_wire214    <= data43x(7 DOWNTO 0);
	sub_wire213    <= data44x(7 DOWNTO 0);
	sub_wire212    <= data45x(7 DOWNTO 0);
	sub_wire211    <= data46x(7 DOWNTO 0);
	sub_wire210    <= data47x(7 DOWNTO 0);
	sub_wire209    <= data48x(7 DOWNTO 0);
	sub_wire208    <= data49x(7 DOWNTO 0);
	sub_wire207    <= data50x(7 DOWNTO 0);
	sub_wire206    <= data51x(7 DOWNTO 0);
	sub_wire205    <= data52x(7 DOWNTO 0);
	sub_wire204    <= data53x(7 DOWNTO 0);
	sub_wire203    <= data54x(7 DOWNTO 0);
	sub_wire202    <= data55x(7 DOWNTO 0);
	sub_wire201    <= data56x(7 DOWNTO 0);
	sub_wire200    <= data57x(7 DOWNTO 0);
	sub_wire199    <= data58x(7 DOWNTO 0);
	sub_wire198    <= data59x(7 DOWNTO 0);
	sub_wire197    <= data60x(7 DOWNTO 0);
	sub_wire196    <= data61x(7 DOWNTO 0);
	sub_wire195    <= data62x(7 DOWNTO 0);
	sub_wire194    <= data63x(7 DOWNTO 0);
	sub_wire193    <= data64x(7 DOWNTO 0);
	sub_wire192    <= data65x(7 DOWNTO 0);
	sub_wire191    <= data66x(7 DOWNTO 0);
	sub_wire190    <= data67x(7 DOWNTO 0);
	sub_wire189    <= data68x(7 DOWNTO 0);
	sub_wire188    <= data69x(7 DOWNTO 0);
	sub_wire187    <= data70x(7 DOWNTO 0);
	sub_wire186    <= data71x(7 DOWNTO 0);
	sub_wire185    <= data72x(7 DOWNTO 0);
	sub_wire184    <= data73x(7 DOWNTO 0);
	sub_wire183    <= data74x(7 DOWNTO 0);
	sub_wire182    <= data75x(7 DOWNTO 0);
	sub_wire181    <= data76x(7 DOWNTO 0);
	sub_wire180    <= data77x(7 DOWNTO 0);
	sub_wire179    <= data78x(7 DOWNTO 0);
	sub_wire178    <= data79x(7 DOWNTO 0);
	sub_wire177    <= data80x(7 DOWNTO 0);
	sub_wire176    <= data81x(7 DOWNTO 0);
	sub_wire175    <= data82x(7 DOWNTO 0);
	sub_wire174    <= data83x(7 DOWNTO 0);
	sub_wire173    <= data84x(7 DOWNTO 0);
	sub_wire172    <= data85x(7 DOWNTO 0);
	sub_wire171    <= data86x(7 DOWNTO 0);
	sub_wire170    <= data87x(7 DOWNTO 0);
	sub_wire169    <= data88x(7 DOWNTO 0);
	sub_wire168    <= data89x(7 DOWNTO 0);
	sub_wire167    <= data90x(7 DOWNTO 0);
	sub_wire166    <= data91x(7 DOWNTO 0);
	sub_wire165    <= data92x(7 DOWNTO 0);
	sub_wire164    <= data93x(7 DOWNTO 0);
	sub_wire163    <= data94x(7 DOWNTO 0);
	sub_wire162    <= data95x(7 DOWNTO 0);
	sub_wire161    <= data96x(7 DOWNTO 0);
	sub_wire160    <= data97x(7 DOWNTO 0);
	sub_wire159    <= data98x(7 DOWNTO 0);
	sub_wire158    <= data99x(7 DOWNTO 0);
	sub_wire157    <= data100x(7 DOWNTO 0);
	sub_wire156    <= data101x(7 DOWNTO 0);
	sub_wire155    <= data102x(7 DOWNTO 0);
	sub_wire154    <= data103x(7 DOWNTO 0);
	sub_wire153    <= data104x(7 DOWNTO 0);
	sub_wire152    <= data105x(7 DOWNTO 0);
	sub_wire151    <= data106x(7 DOWNTO 0);
	sub_wire150    <= data107x(7 DOWNTO 0);
	sub_wire149    <= data108x(7 DOWNTO 0);
	sub_wire148    <= data109x(7 DOWNTO 0);
	sub_wire147    <= data110x(7 DOWNTO 0);
	sub_wire146    <= data111x(7 DOWNTO 0);
	sub_wire145    <= data112x(7 DOWNTO 0);
	sub_wire144    <= data113x(7 DOWNTO 0);
	sub_wire143    <= data114x(7 DOWNTO 0);
	sub_wire142    <= data115x(7 DOWNTO 0);
	sub_wire141    <= data116x(7 DOWNTO 0);
	sub_wire140    <= data117x(7 DOWNTO 0);
	sub_wire139    <= data118x(7 DOWNTO 0);
	sub_wire138    <= data119x(7 DOWNTO 0);
	sub_wire137    <= data120x(7 DOWNTO 0);
	sub_wire136    <= data121x(7 DOWNTO 0);
	sub_wire135    <= data122x(7 DOWNTO 0);
	sub_wire134    <= data123x(7 DOWNTO 0);
	sub_wire133    <= data124x(7 DOWNTO 0);
	sub_wire132    <= data125x(7 DOWNTO 0);
	sub_wire131    <= data126x(7 DOWNTO 0);
	sub_wire130    <= data127x(7 DOWNTO 0);
	sub_wire129    <= data128x(7 DOWNTO 0);
	sub_wire128    <= data129x(7 DOWNTO 0);
	sub_wire127    <= data130x(7 DOWNTO 0);
	sub_wire126    <= data131x(7 DOWNTO 0);
	sub_wire125    <= data132x(7 DOWNTO 0);
	sub_wire124    <= data133x(7 DOWNTO 0);
	sub_wire123    <= data134x(7 DOWNTO 0);
	sub_wire122    <= data135x(7 DOWNTO 0);
	sub_wire121    <= data136x(7 DOWNTO 0);
	sub_wire120    <= data137x(7 DOWNTO 0);
	sub_wire119    <= data138x(7 DOWNTO 0);
	sub_wire118    <= data139x(7 DOWNTO 0);
	sub_wire117    <= data140x(7 DOWNTO 0);
	sub_wire116    <= data141x(7 DOWNTO 0);
	sub_wire115    <= data142x(7 DOWNTO 0);
	sub_wire114    <= data143x(7 DOWNTO 0);
	sub_wire113    <= data144x(7 DOWNTO 0);
	sub_wire112    <= data145x(7 DOWNTO 0);
	sub_wire111    <= data146x(7 DOWNTO 0);
	sub_wire110    <= data147x(7 DOWNTO 0);
	sub_wire109    <= data148x(7 DOWNTO 0);
	sub_wire108    <= data149x(7 DOWNTO 0);
	sub_wire107    <= data150x(7 DOWNTO 0);
	sub_wire106    <= data151x(7 DOWNTO 0);
	sub_wire105    <= data152x(7 DOWNTO 0);
	sub_wire104    <= data153x(7 DOWNTO 0);
	sub_wire103    <= data154x(7 DOWNTO 0);
	sub_wire102    <= data155x(7 DOWNTO 0);
	sub_wire101    <= data156x(7 DOWNTO 0);
	sub_wire100    <= data157x(7 DOWNTO 0);
	sub_wire99    <= data158x(7 DOWNTO 0);
	sub_wire98    <= data159x(7 DOWNTO 0);
	sub_wire97    <= data160x(7 DOWNTO 0);
	sub_wire96    <= data161x(7 DOWNTO 0);
	sub_wire95    <= data162x(7 DOWNTO 0);
	sub_wire94    <= data163x(7 DOWNTO 0);
	sub_wire93    <= data164x(7 DOWNTO 0);
	sub_wire92    <= data165x(7 DOWNTO 0);
	sub_wire91    <= data166x(7 DOWNTO 0);
	sub_wire90    <= data167x(7 DOWNTO 0);
	sub_wire89    <= data168x(7 DOWNTO 0);
	sub_wire88    <= data169x(7 DOWNTO 0);
	sub_wire87    <= data170x(7 DOWNTO 0);
	sub_wire86    <= data171x(7 DOWNTO 0);
	sub_wire85    <= data172x(7 DOWNTO 0);
	sub_wire84    <= data173x(7 DOWNTO 0);
	sub_wire83    <= data174x(7 DOWNTO 0);
	sub_wire82    <= data175x(7 DOWNTO 0);
	sub_wire81    <= data176x(7 DOWNTO 0);
	sub_wire80    <= data177x(7 DOWNTO 0);
	sub_wire79    <= data178x(7 DOWNTO 0);
	sub_wire78    <= data179x(7 DOWNTO 0);
	sub_wire77    <= data180x(7 DOWNTO 0);
	sub_wire76    <= data181x(7 DOWNTO 0);
	sub_wire75    <= data182x(7 DOWNTO 0);
	sub_wire74    <= data183x(7 DOWNTO 0);
	sub_wire73    <= data184x(7 DOWNTO 0);
	sub_wire72    <= data185x(7 DOWNTO 0);
	sub_wire71    <= data186x(7 DOWNTO 0);
	sub_wire70    <= data187x(7 DOWNTO 0);
	sub_wire69    <= data188x(7 DOWNTO 0);
	sub_wire68    <= data189x(7 DOWNTO 0);
	sub_wire67    <= data190x(7 DOWNTO 0);
	sub_wire66    <= data191x(7 DOWNTO 0);
	sub_wire65    <= data192x(7 DOWNTO 0);
	sub_wire64    <= data193x(7 DOWNTO 0);
	sub_wire63    <= data194x(7 DOWNTO 0);
	sub_wire62    <= data195x(7 DOWNTO 0);
	sub_wire61    <= data196x(7 DOWNTO 0);
	sub_wire60    <= data197x(7 DOWNTO 0);
	sub_wire59    <= data198x(7 DOWNTO 0);
	sub_wire58    <= data199x(7 DOWNTO 0);
	sub_wire57    <= data200x(7 DOWNTO 0);
	sub_wire56    <= data201x(7 DOWNTO 0);
	sub_wire55    <= data202x(7 DOWNTO 0);
	sub_wire54    <= data203x(7 DOWNTO 0);
	sub_wire53    <= data204x(7 DOWNTO 0);
	sub_wire52    <= data205x(7 DOWNTO 0);
	sub_wire51    <= data206x(7 DOWNTO 0);
	sub_wire50    <= data207x(7 DOWNTO 0);
	sub_wire49    <= data208x(7 DOWNTO 0);
	sub_wire48    <= data209x(7 DOWNTO 0);
	sub_wire47    <= data210x(7 DOWNTO 0);
	sub_wire46    <= data211x(7 DOWNTO 0);
	sub_wire45    <= data212x(7 DOWNTO 0);
	sub_wire44    <= data213x(7 DOWNTO 0);
	sub_wire43    <= data214x(7 DOWNTO 0);
	sub_wire42    <= data215x(7 DOWNTO 0);
	sub_wire41    <= data216x(7 DOWNTO 0);
	sub_wire40    <= data217x(7 DOWNTO 0);
	sub_wire39    <= data218x(7 DOWNTO 0);
	sub_wire38    <= data219x(7 DOWNTO 0);
	sub_wire37    <= data220x(7 DOWNTO 0);
	sub_wire36    <= data221x(7 DOWNTO 0);
	sub_wire35    <= data222x(7 DOWNTO 0);
	sub_wire34    <= data223x(7 DOWNTO 0);
	sub_wire33    <= data224x(7 DOWNTO 0);
	sub_wire32    <= data225x(7 DOWNTO 0);
	sub_wire31    <= data226x(7 DOWNTO 0);
	sub_wire30    <= data227x(7 DOWNTO 0);
	sub_wire29    <= data228x(7 DOWNTO 0);
	sub_wire28    <= data229x(7 DOWNTO 0);
	sub_wire27    <= data230x(7 DOWNTO 0);
	sub_wire26    <= data231x(7 DOWNTO 0);
	sub_wire25    <= data232x(7 DOWNTO 0);
	sub_wire24    <= data233x(7 DOWNTO 0);
	sub_wire23    <= data234x(7 DOWNTO 0);
	sub_wire22    <= data235x(7 DOWNTO 0);
	sub_wire21    <= data236x(7 DOWNTO 0);
	sub_wire20    <= data237x(7 DOWNTO 0);
	sub_wire19    <= data238x(7 DOWNTO 0);
	sub_wire18    <= data239x(7 DOWNTO 0);
	sub_wire17    <= data240x(7 DOWNTO 0);
	sub_wire16    <= data241x(7 DOWNTO 0);
	sub_wire15    <= data242x(7 DOWNTO 0);
	sub_wire14    <= data243x(7 DOWNTO 0);
	sub_wire13    <= data244x(7 DOWNTO 0);
	sub_wire12    <= data245x(7 DOWNTO 0);
	sub_wire11    <= data246x(7 DOWNTO 0);
	sub_wire10    <= data247x(7 DOWNTO 0);
	sub_wire9    <= data248x(7 DOWNTO 0);
	sub_wire8    <= data249x(7 DOWNTO 0);
	sub_wire7    <= data250x(7 DOWNTO 0);
	sub_wire6    <= data251x(7 DOWNTO 0);
	sub_wire5    <= data252x(7 DOWNTO 0);
	sub_wire4    <= data253x(7 DOWNTO 0);
	sub_wire3    <= data254x(7 DOWNTO 0);
	result    <= sub_wire0(7 DOWNTO 0);
	sub_wire1    <= data255x(7 DOWNTO 0);
	sub_wire2(255, 0)    <= sub_wire1(0);
	sub_wire2(255, 1)    <= sub_wire1(1);
	sub_wire2(255, 2)    <= sub_wire1(2);
	sub_wire2(255, 3)    <= sub_wire1(3);
	sub_wire2(255, 4)    <= sub_wire1(4);
	sub_wire2(255, 5)    <= sub_wire1(5);
	sub_wire2(255, 6)    <= sub_wire1(6);
	sub_wire2(255, 7)    <= sub_wire1(7);
	sub_wire2(254, 0)    <= sub_wire3(0);
	sub_wire2(254, 1)    <= sub_wire3(1);
	sub_wire2(254, 2)    <= sub_wire3(2);
	sub_wire2(254, 3)    <= sub_wire3(3);
	sub_wire2(254, 4)    <= sub_wire3(4);
	sub_wire2(254, 5)    <= sub_wire3(5);
	sub_wire2(254, 6)    <= sub_wire3(6);
	sub_wire2(254, 7)    <= sub_wire3(7);
	sub_wire2(253, 0)    <= sub_wire4(0);
	sub_wire2(253, 1)    <= sub_wire4(1);
	sub_wire2(253, 2)    <= sub_wire4(2);
	sub_wire2(253, 3)    <= sub_wire4(3);
	sub_wire2(253, 4)    <= sub_wire4(4);
	sub_wire2(253, 5)    <= sub_wire4(5);
	sub_wire2(253, 6)    <= sub_wire4(6);
	sub_wire2(253, 7)    <= sub_wire4(7);
	sub_wire2(252, 0)    <= sub_wire5(0);
	sub_wire2(252, 1)    <= sub_wire5(1);
	sub_wire2(252, 2)    <= sub_wire5(2);
	sub_wire2(252, 3)    <= sub_wire5(3);
	sub_wire2(252, 4)    <= sub_wire5(4);
	sub_wire2(252, 5)    <= sub_wire5(5);
	sub_wire2(252, 6)    <= sub_wire5(6);
	sub_wire2(252, 7)    <= sub_wire5(7);
	sub_wire2(251, 0)    <= sub_wire6(0);
	sub_wire2(251, 1)    <= sub_wire6(1);
	sub_wire2(251, 2)    <= sub_wire6(2);
	sub_wire2(251, 3)    <= sub_wire6(3);
	sub_wire2(251, 4)    <= sub_wire6(4);
	sub_wire2(251, 5)    <= sub_wire6(5);
	sub_wire2(251, 6)    <= sub_wire6(6);
	sub_wire2(251, 7)    <= sub_wire6(7);
	sub_wire2(250, 0)    <= sub_wire7(0);
	sub_wire2(250, 1)    <= sub_wire7(1);
	sub_wire2(250, 2)    <= sub_wire7(2);
	sub_wire2(250, 3)    <= sub_wire7(3);
	sub_wire2(250, 4)    <= sub_wire7(4);
	sub_wire2(250, 5)    <= sub_wire7(5);
	sub_wire2(250, 6)    <= sub_wire7(6);
	sub_wire2(250, 7)    <= sub_wire7(7);
	sub_wire2(249, 0)    <= sub_wire8(0);
	sub_wire2(249, 1)    <= sub_wire8(1);
	sub_wire2(249, 2)    <= sub_wire8(2);
	sub_wire2(249, 3)    <= sub_wire8(3);
	sub_wire2(249, 4)    <= sub_wire8(4);
	sub_wire2(249, 5)    <= sub_wire8(5);
	sub_wire2(249, 6)    <= sub_wire8(6);
	sub_wire2(249, 7)    <= sub_wire8(7);
	sub_wire2(248, 0)    <= sub_wire9(0);
	sub_wire2(248, 1)    <= sub_wire9(1);
	sub_wire2(248, 2)    <= sub_wire9(2);
	sub_wire2(248, 3)    <= sub_wire9(3);
	sub_wire2(248, 4)    <= sub_wire9(4);
	sub_wire2(248, 5)    <= sub_wire9(5);
	sub_wire2(248, 6)    <= sub_wire9(6);
	sub_wire2(248, 7)    <= sub_wire9(7);
	sub_wire2(247, 0)    <= sub_wire10(0);
	sub_wire2(247, 1)    <= sub_wire10(1);
	sub_wire2(247, 2)    <= sub_wire10(2);
	sub_wire2(247, 3)    <= sub_wire10(3);
	sub_wire2(247, 4)    <= sub_wire10(4);
	sub_wire2(247, 5)    <= sub_wire10(5);
	sub_wire2(247, 6)    <= sub_wire10(6);
	sub_wire2(247, 7)    <= sub_wire10(7);
	sub_wire2(246, 0)    <= sub_wire11(0);
	sub_wire2(246, 1)    <= sub_wire11(1);
	sub_wire2(246, 2)    <= sub_wire11(2);
	sub_wire2(246, 3)    <= sub_wire11(3);
	sub_wire2(246, 4)    <= sub_wire11(4);
	sub_wire2(246, 5)    <= sub_wire11(5);
	sub_wire2(246, 6)    <= sub_wire11(6);
	sub_wire2(246, 7)    <= sub_wire11(7);
	sub_wire2(245, 0)    <= sub_wire12(0);
	sub_wire2(245, 1)    <= sub_wire12(1);
	sub_wire2(245, 2)    <= sub_wire12(2);
	sub_wire2(245, 3)    <= sub_wire12(3);
	sub_wire2(245, 4)    <= sub_wire12(4);
	sub_wire2(245, 5)    <= sub_wire12(5);
	sub_wire2(245, 6)    <= sub_wire12(6);
	sub_wire2(245, 7)    <= sub_wire12(7);
	sub_wire2(244, 0)    <= sub_wire13(0);
	sub_wire2(244, 1)    <= sub_wire13(1);
	sub_wire2(244, 2)    <= sub_wire13(2);
	sub_wire2(244, 3)    <= sub_wire13(3);
	sub_wire2(244, 4)    <= sub_wire13(4);
	sub_wire2(244, 5)    <= sub_wire13(5);
	sub_wire2(244, 6)    <= sub_wire13(6);
	sub_wire2(244, 7)    <= sub_wire13(7);
	sub_wire2(243, 0)    <= sub_wire14(0);
	sub_wire2(243, 1)    <= sub_wire14(1);
	sub_wire2(243, 2)    <= sub_wire14(2);
	sub_wire2(243, 3)    <= sub_wire14(3);
	sub_wire2(243, 4)    <= sub_wire14(4);
	sub_wire2(243, 5)    <= sub_wire14(5);
	sub_wire2(243, 6)    <= sub_wire14(6);
	sub_wire2(243, 7)    <= sub_wire14(7);
	sub_wire2(242, 0)    <= sub_wire15(0);
	sub_wire2(242, 1)    <= sub_wire15(1);
	sub_wire2(242, 2)    <= sub_wire15(2);
	sub_wire2(242, 3)    <= sub_wire15(3);
	sub_wire2(242, 4)    <= sub_wire15(4);
	sub_wire2(242, 5)    <= sub_wire15(5);
	sub_wire2(242, 6)    <= sub_wire15(6);
	sub_wire2(242, 7)    <= sub_wire15(7);
	sub_wire2(241, 0)    <= sub_wire16(0);
	sub_wire2(241, 1)    <= sub_wire16(1);
	sub_wire2(241, 2)    <= sub_wire16(2);
	sub_wire2(241, 3)    <= sub_wire16(3);
	sub_wire2(241, 4)    <= sub_wire16(4);
	sub_wire2(241, 5)    <= sub_wire16(5);
	sub_wire2(241, 6)    <= sub_wire16(6);
	sub_wire2(241, 7)    <= sub_wire16(7);
	sub_wire2(240, 0)    <= sub_wire17(0);
	sub_wire2(240, 1)    <= sub_wire17(1);
	sub_wire2(240, 2)    <= sub_wire17(2);
	sub_wire2(240, 3)    <= sub_wire17(3);
	sub_wire2(240, 4)    <= sub_wire17(4);
	sub_wire2(240, 5)    <= sub_wire17(5);
	sub_wire2(240, 6)    <= sub_wire17(6);
	sub_wire2(240, 7)    <= sub_wire17(7);
	sub_wire2(239, 0)    <= sub_wire18(0);
	sub_wire2(239, 1)    <= sub_wire18(1);
	sub_wire2(239, 2)    <= sub_wire18(2);
	sub_wire2(239, 3)    <= sub_wire18(3);
	sub_wire2(239, 4)    <= sub_wire18(4);
	sub_wire2(239, 5)    <= sub_wire18(5);
	sub_wire2(239, 6)    <= sub_wire18(6);
	sub_wire2(239, 7)    <= sub_wire18(7);
	sub_wire2(238, 0)    <= sub_wire19(0);
	sub_wire2(238, 1)    <= sub_wire19(1);
	sub_wire2(238, 2)    <= sub_wire19(2);
	sub_wire2(238, 3)    <= sub_wire19(3);
	sub_wire2(238, 4)    <= sub_wire19(4);
	sub_wire2(238, 5)    <= sub_wire19(5);
	sub_wire2(238, 6)    <= sub_wire19(6);
	sub_wire2(238, 7)    <= sub_wire19(7);
	sub_wire2(237, 0)    <= sub_wire20(0);
	sub_wire2(237, 1)    <= sub_wire20(1);
	sub_wire2(237, 2)    <= sub_wire20(2);
	sub_wire2(237, 3)    <= sub_wire20(3);
	sub_wire2(237, 4)    <= sub_wire20(4);
	sub_wire2(237, 5)    <= sub_wire20(5);
	sub_wire2(237, 6)    <= sub_wire20(6);
	sub_wire2(237, 7)    <= sub_wire20(7);
	sub_wire2(236, 0)    <= sub_wire21(0);
	sub_wire2(236, 1)    <= sub_wire21(1);
	sub_wire2(236, 2)    <= sub_wire21(2);
	sub_wire2(236, 3)    <= sub_wire21(3);
	sub_wire2(236, 4)    <= sub_wire21(4);
	sub_wire2(236, 5)    <= sub_wire21(5);
	sub_wire2(236, 6)    <= sub_wire21(6);
	sub_wire2(236, 7)    <= sub_wire21(7);
	sub_wire2(235, 0)    <= sub_wire22(0);
	sub_wire2(235, 1)    <= sub_wire22(1);
	sub_wire2(235, 2)    <= sub_wire22(2);
	sub_wire2(235, 3)    <= sub_wire22(3);
	sub_wire2(235, 4)    <= sub_wire22(4);
	sub_wire2(235, 5)    <= sub_wire22(5);
	sub_wire2(235, 6)    <= sub_wire22(6);
	sub_wire2(235, 7)    <= sub_wire22(7);
	sub_wire2(234, 0)    <= sub_wire23(0);
	sub_wire2(234, 1)    <= sub_wire23(1);
	sub_wire2(234, 2)    <= sub_wire23(2);
	sub_wire2(234, 3)    <= sub_wire23(3);
	sub_wire2(234, 4)    <= sub_wire23(4);
	sub_wire2(234, 5)    <= sub_wire23(5);
	sub_wire2(234, 6)    <= sub_wire23(6);
	sub_wire2(234, 7)    <= sub_wire23(7);
	sub_wire2(233, 0)    <= sub_wire24(0);
	sub_wire2(233, 1)    <= sub_wire24(1);
	sub_wire2(233, 2)    <= sub_wire24(2);
	sub_wire2(233, 3)    <= sub_wire24(3);
	sub_wire2(233, 4)    <= sub_wire24(4);
	sub_wire2(233, 5)    <= sub_wire24(5);
	sub_wire2(233, 6)    <= sub_wire24(6);
	sub_wire2(233, 7)    <= sub_wire24(7);
	sub_wire2(232, 0)    <= sub_wire25(0);
	sub_wire2(232, 1)    <= sub_wire25(1);
	sub_wire2(232, 2)    <= sub_wire25(2);
	sub_wire2(232, 3)    <= sub_wire25(3);
	sub_wire2(232, 4)    <= sub_wire25(4);
	sub_wire2(232, 5)    <= sub_wire25(5);
	sub_wire2(232, 6)    <= sub_wire25(6);
	sub_wire2(232, 7)    <= sub_wire25(7);
	sub_wire2(231, 0)    <= sub_wire26(0);
	sub_wire2(231, 1)    <= sub_wire26(1);
	sub_wire2(231, 2)    <= sub_wire26(2);
	sub_wire2(231, 3)    <= sub_wire26(3);
	sub_wire2(231, 4)    <= sub_wire26(4);
	sub_wire2(231, 5)    <= sub_wire26(5);
	sub_wire2(231, 6)    <= sub_wire26(6);
	sub_wire2(231, 7)    <= sub_wire26(7);
	sub_wire2(230, 0)    <= sub_wire27(0);
	sub_wire2(230, 1)    <= sub_wire27(1);
	sub_wire2(230, 2)    <= sub_wire27(2);
	sub_wire2(230, 3)    <= sub_wire27(3);
	sub_wire2(230, 4)    <= sub_wire27(4);
	sub_wire2(230, 5)    <= sub_wire27(5);
	sub_wire2(230, 6)    <= sub_wire27(6);
	sub_wire2(230, 7)    <= sub_wire27(7);
	sub_wire2(229, 0)    <= sub_wire28(0);
	sub_wire2(229, 1)    <= sub_wire28(1);
	sub_wire2(229, 2)    <= sub_wire28(2);
	sub_wire2(229, 3)    <= sub_wire28(3);
	sub_wire2(229, 4)    <= sub_wire28(4);
	sub_wire2(229, 5)    <= sub_wire28(5);
	sub_wire2(229, 6)    <= sub_wire28(6);
	sub_wire2(229, 7)    <= sub_wire28(7);
	sub_wire2(228, 0)    <= sub_wire29(0);
	sub_wire2(228, 1)    <= sub_wire29(1);
	sub_wire2(228, 2)    <= sub_wire29(2);
	sub_wire2(228, 3)    <= sub_wire29(3);
	sub_wire2(228, 4)    <= sub_wire29(4);
	sub_wire2(228, 5)    <= sub_wire29(5);
	sub_wire2(228, 6)    <= sub_wire29(6);
	sub_wire2(228, 7)    <= sub_wire29(7);
	sub_wire2(227, 0)    <= sub_wire30(0);
	sub_wire2(227, 1)    <= sub_wire30(1);
	sub_wire2(227, 2)    <= sub_wire30(2);
	sub_wire2(227, 3)    <= sub_wire30(3);
	sub_wire2(227, 4)    <= sub_wire30(4);
	sub_wire2(227, 5)    <= sub_wire30(5);
	sub_wire2(227, 6)    <= sub_wire30(6);
	sub_wire2(227, 7)    <= sub_wire30(7);
	sub_wire2(226, 0)    <= sub_wire31(0);
	sub_wire2(226, 1)    <= sub_wire31(1);
	sub_wire2(226, 2)    <= sub_wire31(2);
	sub_wire2(226, 3)    <= sub_wire31(3);
	sub_wire2(226, 4)    <= sub_wire31(4);
	sub_wire2(226, 5)    <= sub_wire31(5);
	sub_wire2(226, 6)    <= sub_wire31(6);
	sub_wire2(226, 7)    <= sub_wire31(7);
	sub_wire2(225, 0)    <= sub_wire32(0);
	sub_wire2(225, 1)    <= sub_wire32(1);
	sub_wire2(225, 2)    <= sub_wire32(2);
	sub_wire2(225, 3)    <= sub_wire32(3);
	sub_wire2(225, 4)    <= sub_wire32(4);
	sub_wire2(225, 5)    <= sub_wire32(5);
	sub_wire2(225, 6)    <= sub_wire32(6);
	sub_wire2(225, 7)    <= sub_wire32(7);
	sub_wire2(224, 0)    <= sub_wire33(0);
	sub_wire2(224, 1)    <= sub_wire33(1);
	sub_wire2(224, 2)    <= sub_wire33(2);
	sub_wire2(224, 3)    <= sub_wire33(3);
	sub_wire2(224, 4)    <= sub_wire33(4);
	sub_wire2(224, 5)    <= sub_wire33(5);
	sub_wire2(224, 6)    <= sub_wire33(6);
	sub_wire2(224, 7)    <= sub_wire33(7);
	sub_wire2(223, 0)    <= sub_wire34(0);
	sub_wire2(223, 1)    <= sub_wire34(1);
	sub_wire2(223, 2)    <= sub_wire34(2);
	sub_wire2(223, 3)    <= sub_wire34(3);
	sub_wire2(223, 4)    <= sub_wire34(4);
	sub_wire2(223, 5)    <= sub_wire34(5);
	sub_wire2(223, 6)    <= sub_wire34(6);
	sub_wire2(223, 7)    <= sub_wire34(7);
	sub_wire2(222, 0)    <= sub_wire35(0);
	sub_wire2(222, 1)    <= sub_wire35(1);
	sub_wire2(222, 2)    <= sub_wire35(2);
	sub_wire2(222, 3)    <= sub_wire35(3);
	sub_wire2(222, 4)    <= sub_wire35(4);
	sub_wire2(222, 5)    <= sub_wire35(5);
	sub_wire2(222, 6)    <= sub_wire35(6);
	sub_wire2(222, 7)    <= sub_wire35(7);
	sub_wire2(221, 0)    <= sub_wire36(0);
	sub_wire2(221, 1)    <= sub_wire36(1);
	sub_wire2(221, 2)    <= sub_wire36(2);
	sub_wire2(221, 3)    <= sub_wire36(3);
	sub_wire2(221, 4)    <= sub_wire36(4);
	sub_wire2(221, 5)    <= sub_wire36(5);
	sub_wire2(221, 6)    <= sub_wire36(6);
	sub_wire2(221, 7)    <= sub_wire36(7);
	sub_wire2(220, 0)    <= sub_wire37(0);
	sub_wire2(220, 1)    <= sub_wire37(1);
	sub_wire2(220, 2)    <= sub_wire37(2);
	sub_wire2(220, 3)    <= sub_wire37(3);
	sub_wire2(220, 4)    <= sub_wire37(4);
	sub_wire2(220, 5)    <= sub_wire37(5);
	sub_wire2(220, 6)    <= sub_wire37(6);
	sub_wire2(220, 7)    <= sub_wire37(7);
	sub_wire2(219, 0)    <= sub_wire38(0);
	sub_wire2(219, 1)    <= sub_wire38(1);
	sub_wire2(219, 2)    <= sub_wire38(2);
	sub_wire2(219, 3)    <= sub_wire38(3);
	sub_wire2(219, 4)    <= sub_wire38(4);
	sub_wire2(219, 5)    <= sub_wire38(5);
	sub_wire2(219, 6)    <= sub_wire38(6);
	sub_wire2(219, 7)    <= sub_wire38(7);
	sub_wire2(218, 0)    <= sub_wire39(0);
	sub_wire2(218, 1)    <= sub_wire39(1);
	sub_wire2(218, 2)    <= sub_wire39(2);
	sub_wire2(218, 3)    <= sub_wire39(3);
	sub_wire2(218, 4)    <= sub_wire39(4);
	sub_wire2(218, 5)    <= sub_wire39(5);
	sub_wire2(218, 6)    <= sub_wire39(6);
	sub_wire2(218, 7)    <= sub_wire39(7);
	sub_wire2(217, 0)    <= sub_wire40(0);
	sub_wire2(217, 1)    <= sub_wire40(1);
	sub_wire2(217, 2)    <= sub_wire40(2);
	sub_wire2(217, 3)    <= sub_wire40(3);
	sub_wire2(217, 4)    <= sub_wire40(4);
	sub_wire2(217, 5)    <= sub_wire40(5);
	sub_wire2(217, 6)    <= sub_wire40(6);
	sub_wire2(217, 7)    <= sub_wire40(7);
	sub_wire2(216, 0)    <= sub_wire41(0);
	sub_wire2(216, 1)    <= sub_wire41(1);
	sub_wire2(216, 2)    <= sub_wire41(2);
	sub_wire2(216, 3)    <= sub_wire41(3);
	sub_wire2(216, 4)    <= sub_wire41(4);
	sub_wire2(216, 5)    <= sub_wire41(5);
	sub_wire2(216, 6)    <= sub_wire41(6);
	sub_wire2(216, 7)    <= sub_wire41(7);
	sub_wire2(215, 0)    <= sub_wire42(0);
	sub_wire2(215, 1)    <= sub_wire42(1);
	sub_wire2(215, 2)    <= sub_wire42(2);
	sub_wire2(215, 3)    <= sub_wire42(3);
	sub_wire2(215, 4)    <= sub_wire42(4);
	sub_wire2(215, 5)    <= sub_wire42(5);
	sub_wire2(215, 6)    <= sub_wire42(6);
	sub_wire2(215, 7)    <= sub_wire42(7);
	sub_wire2(214, 0)    <= sub_wire43(0);
	sub_wire2(214, 1)    <= sub_wire43(1);
	sub_wire2(214, 2)    <= sub_wire43(2);
	sub_wire2(214, 3)    <= sub_wire43(3);
	sub_wire2(214, 4)    <= sub_wire43(4);
	sub_wire2(214, 5)    <= sub_wire43(5);
	sub_wire2(214, 6)    <= sub_wire43(6);
	sub_wire2(214, 7)    <= sub_wire43(7);
	sub_wire2(213, 0)    <= sub_wire44(0);
	sub_wire2(213, 1)    <= sub_wire44(1);
	sub_wire2(213, 2)    <= sub_wire44(2);
	sub_wire2(213, 3)    <= sub_wire44(3);
	sub_wire2(213, 4)    <= sub_wire44(4);
	sub_wire2(213, 5)    <= sub_wire44(5);
	sub_wire2(213, 6)    <= sub_wire44(6);
	sub_wire2(213, 7)    <= sub_wire44(7);
	sub_wire2(212, 0)    <= sub_wire45(0);
	sub_wire2(212, 1)    <= sub_wire45(1);
	sub_wire2(212, 2)    <= sub_wire45(2);
	sub_wire2(212, 3)    <= sub_wire45(3);
	sub_wire2(212, 4)    <= sub_wire45(4);
	sub_wire2(212, 5)    <= sub_wire45(5);
	sub_wire2(212, 6)    <= sub_wire45(6);
	sub_wire2(212, 7)    <= sub_wire45(7);
	sub_wire2(211, 0)    <= sub_wire46(0);
	sub_wire2(211, 1)    <= sub_wire46(1);
	sub_wire2(211, 2)    <= sub_wire46(2);
	sub_wire2(211, 3)    <= sub_wire46(3);
	sub_wire2(211, 4)    <= sub_wire46(4);
	sub_wire2(211, 5)    <= sub_wire46(5);
	sub_wire2(211, 6)    <= sub_wire46(6);
	sub_wire2(211, 7)    <= sub_wire46(7);
	sub_wire2(210, 0)    <= sub_wire47(0);
	sub_wire2(210, 1)    <= sub_wire47(1);
	sub_wire2(210, 2)    <= sub_wire47(2);
	sub_wire2(210, 3)    <= sub_wire47(3);
	sub_wire2(210, 4)    <= sub_wire47(4);
	sub_wire2(210, 5)    <= sub_wire47(5);
	sub_wire2(210, 6)    <= sub_wire47(6);
	sub_wire2(210, 7)    <= sub_wire47(7);
	sub_wire2(209, 0)    <= sub_wire48(0);
	sub_wire2(209, 1)    <= sub_wire48(1);
	sub_wire2(209, 2)    <= sub_wire48(2);
	sub_wire2(209, 3)    <= sub_wire48(3);
	sub_wire2(209, 4)    <= sub_wire48(4);
	sub_wire2(209, 5)    <= sub_wire48(5);
	sub_wire2(209, 6)    <= sub_wire48(6);
	sub_wire2(209, 7)    <= sub_wire48(7);
	sub_wire2(208, 0)    <= sub_wire49(0);
	sub_wire2(208, 1)    <= sub_wire49(1);
	sub_wire2(208, 2)    <= sub_wire49(2);
	sub_wire2(208, 3)    <= sub_wire49(3);
	sub_wire2(208, 4)    <= sub_wire49(4);
	sub_wire2(208, 5)    <= sub_wire49(5);
	sub_wire2(208, 6)    <= sub_wire49(6);
	sub_wire2(208, 7)    <= sub_wire49(7);
	sub_wire2(207, 0)    <= sub_wire50(0);
	sub_wire2(207, 1)    <= sub_wire50(1);
	sub_wire2(207, 2)    <= sub_wire50(2);
	sub_wire2(207, 3)    <= sub_wire50(3);
	sub_wire2(207, 4)    <= sub_wire50(4);
	sub_wire2(207, 5)    <= sub_wire50(5);
	sub_wire2(207, 6)    <= sub_wire50(6);
	sub_wire2(207, 7)    <= sub_wire50(7);
	sub_wire2(206, 0)    <= sub_wire51(0);
	sub_wire2(206, 1)    <= sub_wire51(1);
	sub_wire2(206, 2)    <= sub_wire51(2);
	sub_wire2(206, 3)    <= sub_wire51(3);
	sub_wire2(206, 4)    <= sub_wire51(4);
	sub_wire2(206, 5)    <= sub_wire51(5);
	sub_wire2(206, 6)    <= sub_wire51(6);
	sub_wire2(206, 7)    <= sub_wire51(7);
	sub_wire2(205, 0)    <= sub_wire52(0);
	sub_wire2(205, 1)    <= sub_wire52(1);
	sub_wire2(205, 2)    <= sub_wire52(2);
	sub_wire2(205, 3)    <= sub_wire52(3);
	sub_wire2(205, 4)    <= sub_wire52(4);
	sub_wire2(205, 5)    <= sub_wire52(5);
	sub_wire2(205, 6)    <= sub_wire52(6);
	sub_wire2(205, 7)    <= sub_wire52(7);
	sub_wire2(204, 0)    <= sub_wire53(0);
	sub_wire2(204, 1)    <= sub_wire53(1);
	sub_wire2(204, 2)    <= sub_wire53(2);
	sub_wire2(204, 3)    <= sub_wire53(3);
	sub_wire2(204, 4)    <= sub_wire53(4);
	sub_wire2(204, 5)    <= sub_wire53(5);
	sub_wire2(204, 6)    <= sub_wire53(6);
	sub_wire2(204, 7)    <= sub_wire53(7);
	sub_wire2(203, 0)    <= sub_wire54(0);
	sub_wire2(203, 1)    <= sub_wire54(1);
	sub_wire2(203, 2)    <= sub_wire54(2);
	sub_wire2(203, 3)    <= sub_wire54(3);
	sub_wire2(203, 4)    <= sub_wire54(4);
	sub_wire2(203, 5)    <= sub_wire54(5);
	sub_wire2(203, 6)    <= sub_wire54(6);
	sub_wire2(203, 7)    <= sub_wire54(7);
	sub_wire2(202, 0)    <= sub_wire55(0);
	sub_wire2(202, 1)    <= sub_wire55(1);
	sub_wire2(202, 2)    <= sub_wire55(2);
	sub_wire2(202, 3)    <= sub_wire55(3);
	sub_wire2(202, 4)    <= sub_wire55(4);
	sub_wire2(202, 5)    <= sub_wire55(5);
	sub_wire2(202, 6)    <= sub_wire55(6);
	sub_wire2(202, 7)    <= sub_wire55(7);
	sub_wire2(201, 0)    <= sub_wire56(0);
	sub_wire2(201, 1)    <= sub_wire56(1);
	sub_wire2(201, 2)    <= sub_wire56(2);
	sub_wire2(201, 3)    <= sub_wire56(3);
	sub_wire2(201, 4)    <= sub_wire56(4);
	sub_wire2(201, 5)    <= sub_wire56(5);
	sub_wire2(201, 6)    <= sub_wire56(6);
	sub_wire2(201, 7)    <= sub_wire56(7);
	sub_wire2(200, 0)    <= sub_wire57(0);
	sub_wire2(200, 1)    <= sub_wire57(1);
	sub_wire2(200, 2)    <= sub_wire57(2);
	sub_wire2(200, 3)    <= sub_wire57(3);
	sub_wire2(200, 4)    <= sub_wire57(4);
	sub_wire2(200, 5)    <= sub_wire57(5);
	sub_wire2(200, 6)    <= sub_wire57(6);
	sub_wire2(200, 7)    <= sub_wire57(7);
	sub_wire2(199, 0)    <= sub_wire58(0);
	sub_wire2(199, 1)    <= sub_wire58(1);
	sub_wire2(199, 2)    <= sub_wire58(2);
	sub_wire2(199, 3)    <= sub_wire58(3);
	sub_wire2(199, 4)    <= sub_wire58(4);
	sub_wire2(199, 5)    <= sub_wire58(5);
	sub_wire2(199, 6)    <= sub_wire58(6);
	sub_wire2(199, 7)    <= sub_wire58(7);
	sub_wire2(198, 0)    <= sub_wire59(0);
	sub_wire2(198, 1)    <= sub_wire59(1);
	sub_wire2(198, 2)    <= sub_wire59(2);
	sub_wire2(198, 3)    <= sub_wire59(3);
	sub_wire2(198, 4)    <= sub_wire59(4);
	sub_wire2(198, 5)    <= sub_wire59(5);
	sub_wire2(198, 6)    <= sub_wire59(6);
	sub_wire2(198, 7)    <= sub_wire59(7);
	sub_wire2(197, 0)    <= sub_wire60(0);
	sub_wire2(197, 1)    <= sub_wire60(1);
	sub_wire2(197, 2)    <= sub_wire60(2);
	sub_wire2(197, 3)    <= sub_wire60(3);
	sub_wire2(197, 4)    <= sub_wire60(4);
	sub_wire2(197, 5)    <= sub_wire60(5);
	sub_wire2(197, 6)    <= sub_wire60(6);
	sub_wire2(197, 7)    <= sub_wire60(7);
	sub_wire2(196, 0)    <= sub_wire61(0);
	sub_wire2(196, 1)    <= sub_wire61(1);
	sub_wire2(196, 2)    <= sub_wire61(2);
	sub_wire2(196, 3)    <= sub_wire61(3);
	sub_wire2(196, 4)    <= sub_wire61(4);
	sub_wire2(196, 5)    <= sub_wire61(5);
	sub_wire2(196, 6)    <= sub_wire61(6);
	sub_wire2(196, 7)    <= sub_wire61(7);
	sub_wire2(195, 0)    <= sub_wire62(0);
	sub_wire2(195, 1)    <= sub_wire62(1);
	sub_wire2(195, 2)    <= sub_wire62(2);
	sub_wire2(195, 3)    <= sub_wire62(3);
	sub_wire2(195, 4)    <= sub_wire62(4);
	sub_wire2(195, 5)    <= sub_wire62(5);
	sub_wire2(195, 6)    <= sub_wire62(6);
	sub_wire2(195, 7)    <= sub_wire62(7);
	sub_wire2(194, 0)    <= sub_wire63(0);
	sub_wire2(194, 1)    <= sub_wire63(1);
	sub_wire2(194, 2)    <= sub_wire63(2);
	sub_wire2(194, 3)    <= sub_wire63(3);
	sub_wire2(194, 4)    <= sub_wire63(4);
	sub_wire2(194, 5)    <= sub_wire63(5);
	sub_wire2(194, 6)    <= sub_wire63(6);
	sub_wire2(194, 7)    <= sub_wire63(7);
	sub_wire2(193, 0)    <= sub_wire64(0);
	sub_wire2(193, 1)    <= sub_wire64(1);
	sub_wire2(193, 2)    <= sub_wire64(2);
	sub_wire2(193, 3)    <= sub_wire64(3);
	sub_wire2(193, 4)    <= sub_wire64(4);
	sub_wire2(193, 5)    <= sub_wire64(5);
	sub_wire2(193, 6)    <= sub_wire64(6);
	sub_wire2(193, 7)    <= sub_wire64(7);
	sub_wire2(192, 0)    <= sub_wire65(0);
	sub_wire2(192, 1)    <= sub_wire65(1);
	sub_wire2(192, 2)    <= sub_wire65(2);
	sub_wire2(192, 3)    <= sub_wire65(3);
	sub_wire2(192, 4)    <= sub_wire65(4);
	sub_wire2(192, 5)    <= sub_wire65(5);
	sub_wire2(192, 6)    <= sub_wire65(6);
	sub_wire2(192, 7)    <= sub_wire65(7);
	sub_wire2(191, 0)    <= sub_wire66(0);
	sub_wire2(191, 1)    <= sub_wire66(1);
	sub_wire2(191, 2)    <= sub_wire66(2);
	sub_wire2(191, 3)    <= sub_wire66(3);
	sub_wire2(191, 4)    <= sub_wire66(4);
	sub_wire2(191, 5)    <= sub_wire66(5);
	sub_wire2(191, 6)    <= sub_wire66(6);
	sub_wire2(191, 7)    <= sub_wire66(7);
	sub_wire2(190, 0)    <= sub_wire67(0);
	sub_wire2(190, 1)    <= sub_wire67(1);
	sub_wire2(190, 2)    <= sub_wire67(2);
	sub_wire2(190, 3)    <= sub_wire67(3);
	sub_wire2(190, 4)    <= sub_wire67(4);
	sub_wire2(190, 5)    <= sub_wire67(5);
	sub_wire2(190, 6)    <= sub_wire67(6);
	sub_wire2(190, 7)    <= sub_wire67(7);
	sub_wire2(189, 0)    <= sub_wire68(0);
	sub_wire2(189, 1)    <= sub_wire68(1);
	sub_wire2(189, 2)    <= sub_wire68(2);
	sub_wire2(189, 3)    <= sub_wire68(3);
	sub_wire2(189, 4)    <= sub_wire68(4);
	sub_wire2(189, 5)    <= sub_wire68(5);
	sub_wire2(189, 6)    <= sub_wire68(6);
	sub_wire2(189, 7)    <= sub_wire68(7);
	sub_wire2(188, 0)    <= sub_wire69(0);
	sub_wire2(188, 1)    <= sub_wire69(1);
	sub_wire2(188, 2)    <= sub_wire69(2);
	sub_wire2(188, 3)    <= sub_wire69(3);
	sub_wire2(188, 4)    <= sub_wire69(4);
	sub_wire2(188, 5)    <= sub_wire69(5);
	sub_wire2(188, 6)    <= sub_wire69(6);
	sub_wire2(188, 7)    <= sub_wire69(7);
	sub_wire2(187, 0)    <= sub_wire70(0);
	sub_wire2(187, 1)    <= sub_wire70(1);
	sub_wire2(187, 2)    <= sub_wire70(2);
	sub_wire2(187, 3)    <= sub_wire70(3);
	sub_wire2(187, 4)    <= sub_wire70(4);
	sub_wire2(187, 5)    <= sub_wire70(5);
	sub_wire2(187, 6)    <= sub_wire70(6);
	sub_wire2(187, 7)    <= sub_wire70(7);
	sub_wire2(186, 0)    <= sub_wire71(0);
	sub_wire2(186, 1)    <= sub_wire71(1);
	sub_wire2(186, 2)    <= sub_wire71(2);
	sub_wire2(186, 3)    <= sub_wire71(3);
	sub_wire2(186, 4)    <= sub_wire71(4);
	sub_wire2(186, 5)    <= sub_wire71(5);
	sub_wire2(186, 6)    <= sub_wire71(6);
	sub_wire2(186, 7)    <= sub_wire71(7);
	sub_wire2(185, 0)    <= sub_wire72(0);
	sub_wire2(185, 1)    <= sub_wire72(1);
	sub_wire2(185, 2)    <= sub_wire72(2);
	sub_wire2(185, 3)    <= sub_wire72(3);
	sub_wire2(185, 4)    <= sub_wire72(4);
	sub_wire2(185, 5)    <= sub_wire72(5);
	sub_wire2(185, 6)    <= sub_wire72(6);
	sub_wire2(185, 7)    <= sub_wire72(7);
	sub_wire2(184, 0)    <= sub_wire73(0);
	sub_wire2(184, 1)    <= sub_wire73(1);
	sub_wire2(184, 2)    <= sub_wire73(2);
	sub_wire2(184, 3)    <= sub_wire73(3);
	sub_wire2(184, 4)    <= sub_wire73(4);
	sub_wire2(184, 5)    <= sub_wire73(5);
	sub_wire2(184, 6)    <= sub_wire73(6);
	sub_wire2(184, 7)    <= sub_wire73(7);
	sub_wire2(183, 0)    <= sub_wire74(0);
	sub_wire2(183, 1)    <= sub_wire74(1);
	sub_wire2(183, 2)    <= sub_wire74(2);
	sub_wire2(183, 3)    <= sub_wire74(3);
	sub_wire2(183, 4)    <= sub_wire74(4);
	sub_wire2(183, 5)    <= sub_wire74(5);
	sub_wire2(183, 6)    <= sub_wire74(6);
	sub_wire2(183, 7)    <= sub_wire74(7);
	sub_wire2(182, 0)    <= sub_wire75(0);
	sub_wire2(182, 1)    <= sub_wire75(1);
	sub_wire2(182, 2)    <= sub_wire75(2);
	sub_wire2(182, 3)    <= sub_wire75(3);
	sub_wire2(182, 4)    <= sub_wire75(4);
	sub_wire2(182, 5)    <= sub_wire75(5);
	sub_wire2(182, 6)    <= sub_wire75(6);
	sub_wire2(182, 7)    <= sub_wire75(7);
	sub_wire2(181, 0)    <= sub_wire76(0);
	sub_wire2(181, 1)    <= sub_wire76(1);
	sub_wire2(181, 2)    <= sub_wire76(2);
	sub_wire2(181, 3)    <= sub_wire76(3);
	sub_wire2(181, 4)    <= sub_wire76(4);
	sub_wire2(181, 5)    <= sub_wire76(5);
	sub_wire2(181, 6)    <= sub_wire76(6);
	sub_wire2(181, 7)    <= sub_wire76(7);
	sub_wire2(180, 0)    <= sub_wire77(0);
	sub_wire2(180, 1)    <= sub_wire77(1);
	sub_wire2(180, 2)    <= sub_wire77(2);
	sub_wire2(180, 3)    <= sub_wire77(3);
	sub_wire2(180, 4)    <= sub_wire77(4);
	sub_wire2(180, 5)    <= sub_wire77(5);
	sub_wire2(180, 6)    <= sub_wire77(6);
	sub_wire2(180, 7)    <= sub_wire77(7);
	sub_wire2(179, 0)    <= sub_wire78(0);
	sub_wire2(179, 1)    <= sub_wire78(1);
	sub_wire2(179, 2)    <= sub_wire78(2);
	sub_wire2(179, 3)    <= sub_wire78(3);
	sub_wire2(179, 4)    <= sub_wire78(4);
	sub_wire2(179, 5)    <= sub_wire78(5);
	sub_wire2(179, 6)    <= sub_wire78(6);
	sub_wire2(179, 7)    <= sub_wire78(7);
	sub_wire2(178, 0)    <= sub_wire79(0);
	sub_wire2(178, 1)    <= sub_wire79(1);
	sub_wire2(178, 2)    <= sub_wire79(2);
	sub_wire2(178, 3)    <= sub_wire79(3);
	sub_wire2(178, 4)    <= sub_wire79(4);
	sub_wire2(178, 5)    <= sub_wire79(5);
	sub_wire2(178, 6)    <= sub_wire79(6);
	sub_wire2(178, 7)    <= sub_wire79(7);
	sub_wire2(177, 0)    <= sub_wire80(0);
	sub_wire2(177, 1)    <= sub_wire80(1);
	sub_wire2(177, 2)    <= sub_wire80(2);
	sub_wire2(177, 3)    <= sub_wire80(3);
	sub_wire2(177, 4)    <= sub_wire80(4);
	sub_wire2(177, 5)    <= sub_wire80(5);
	sub_wire2(177, 6)    <= sub_wire80(6);
	sub_wire2(177, 7)    <= sub_wire80(7);
	sub_wire2(176, 0)    <= sub_wire81(0);
	sub_wire2(176, 1)    <= sub_wire81(1);
	sub_wire2(176, 2)    <= sub_wire81(2);
	sub_wire2(176, 3)    <= sub_wire81(3);
	sub_wire2(176, 4)    <= sub_wire81(4);
	sub_wire2(176, 5)    <= sub_wire81(5);
	sub_wire2(176, 6)    <= sub_wire81(6);
	sub_wire2(176, 7)    <= sub_wire81(7);
	sub_wire2(175, 0)    <= sub_wire82(0);
	sub_wire2(175, 1)    <= sub_wire82(1);
	sub_wire2(175, 2)    <= sub_wire82(2);
	sub_wire2(175, 3)    <= sub_wire82(3);
	sub_wire2(175, 4)    <= sub_wire82(4);
	sub_wire2(175, 5)    <= sub_wire82(5);
	sub_wire2(175, 6)    <= sub_wire82(6);
	sub_wire2(175, 7)    <= sub_wire82(7);
	sub_wire2(174, 0)    <= sub_wire83(0);
	sub_wire2(174, 1)    <= sub_wire83(1);
	sub_wire2(174, 2)    <= sub_wire83(2);
	sub_wire2(174, 3)    <= sub_wire83(3);
	sub_wire2(174, 4)    <= sub_wire83(4);
	sub_wire2(174, 5)    <= sub_wire83(5);
	sub_wire2(174, 6)    <= sub_wire83(6);
	sub_wire2(174, 7)    <= sub_wire83(7);
	sub_wire2(173, 0)    <= sub_wire84(0);
	sub_wire2(173, 1)    <= sub_wire84(1);
	sub_wire2(173, 2)    <= sub_wire84(2);
	sub_wire2(173, 3)    <= sub_wire84(3);
	sub_wire2(173, 4)    <= sub_wire84(4);
	sub_wire2(173, 5)    <= sub_wire84(5);
	sub_wire2(173, 6)    <= sub_wire84(6);
	sub_wire2(173, 7)    <= sub_wire84(7);
	sub_wire2(172, 0)    <= sub_wire85(0);
	sub_wire2(172, 1)    <= sub_wire85(1);
	sub_wire2(172, 2)    <= sub_wire85(2);
	sub_wire2(172, 3)    <= sub_wire85(3);
	sub_wire2(172, 4)    <= sub_wire85(4);
	sub_wire2(172, 5)    <= sub_wire85(5);
	sub_wire2(172, 6)    <= sub_wire85(6);
	sub_wire2(172, 7)    <= sub_wire85(7);
	sub_wire2(171, 0)    <= sub_wire86(0);
	sub_wire2(171, 1)    <= sub_wire86(1);
	sub_wire2(171, 2)    <= sub_wire86(2);
	sub_wire2(171, 3)    <= sub_wire86(3);
	sub_wire2(171, 4)    <= sub_wire86(4);
	sub_wire2(171, 5)    <= sub_wire86(5);
	sub_wire2(171, 6)    <= sub_wire86(6);
	sub_wire2(171, 7)    <= sub_wire86(7);
	sub_wire2(170, 0)    <= sub_wire87(0);
	sub_wire2(170, 1)    <= sub_wire87(1);
	sub_wire2(170, 2)    <= sub_wire87(2);
	sub_wire2(170, 3)    <= sub_wire87(3);
	sub_wire2(170, 4)    <= sub_wire87(4);
	sub_wire2(170, 5)    <= sub_wire87(5);
	sub_wire2(170, 6)    <= sub_wire87(6);
	sub_wire2(170, 7)    <= sub_wire87(7);
	sub_wire2(169, 0)    <= sub_wire88(0);
	sub_wire2(169, 1)    <= sub_wire88(1);
	sub_wire2(169, 2)    <= sub_wire88(2);
	sub_wire2(169, 3)    <= sub_wire88(3);
	sub_wire2(169, 4)    <= sub_wire88(4);
	sub_wire2(169, 5)    <= sub_wire88(5);
	sub_wire2(169, 6)    <= sub_wire88(6);
	sub_wire2(169, 7)    <= sub_wire88(7);
	sub_wire2(168, 0)    <= sub_wire89(0);
	sub_wire2(168, 1)    <= sub_wire89(1);
	sub_wire2(168, 2)    <= sub_wire89(2);
	sub_wire2(168, 3)    <= sub_wire89(3);
	sub_wire2(168, 4)    <= sub_wire89(4);
	sub_wire2(168, 5)    <= sub_wire89(5);
	sub_wire2(168, 6)    <= sub_wire89(6);
	sub_wire2(168, 7)    <= sub_wire89(7);
	sub_wire2(167, 0)    <= sub_wire90(0);
	sub_wire2(167, 1)    <= sub_wire90(1);
	sub_wire2(167, 2)    <= sub_wire90(2);
	sub_wire2(167, 3)    <= sub_wire90(3);
	sub_wire2(167, 4)    <= sub_wire90(4);
	sub_wire2(167, 5)    <= sub_wire90(5);
	sub_wire2(167, 6)    <= sub_wire90(6);
	sub_wire2(167, 7)    <= sub_wire90(7);
	sub_wire2(166, 0)    <= sub_wire91(0);
	sub_wire2(166, 1)    <= sub_wire91(1);
	sub_wire2(166, 2)    <= sub_wire91(2);
	sub_wire2(166, 3)    <= sub_wire91(3);
	sub_wire2(166, 4)    <= sub_wire91(4);
	sub_wire2(166, 5)    <= sub_wire91(5);
	sub_wire2(166, 6)    <= sub_wire91(6);
	sub_wire2(166, 7)    <= sub_wire91(7);
	sub_wire2(165, 0)    <= sub_wire92(0);
	sub_wire2(165, 1)    <= sub_wire92(1);
	sub_wire2(165, 2)    <= sub_wire92(2);
	sub_wire2(165, 3)    <= sub_wire92(3);
	sub_wire2(165, 4)    <= sub_wire92(4);
	sub_wire2(165, 5)    <= sub_wire92(5);
	sub_wire2(165, 6)    <= sub_wire92(6);
	sub_wire2(165, 7)    <= sub_wire92(7);
	sub_wire2(164, 0)    <= sub_wire93(0);
	sub_wire2(164, 1)    <= sub_wire93(1);
	sub_wire2(164, 2)    <= sub_wire93(2);
	sub_wire2(164, 3)    <= sub_wire93(3);
	sub_wire2(164, 4)    <= sub_wire93(4);
	sub_wire2(164, 5)    <= sub_wire93(5);
	sub_wire2(164, 6)    <= sub_wire93(6);
	sub_wire2(164, 7)    <= sub_wire93(7);
	sub_wire2(163, 0)    <= sub_wire94(0);
	sub_wire2(163, 1)    <= sub_wire94(1);
	sub_wire2(163, 2)    <= sub_wire94(2);
	sub_wire2(163, 3)    <= sub_wire94(3);
	sub_wire2(163, 4)    <= sub_wire94(4);
	sub_wire2(163, 5)    <= sub_wire94(5);
	sub_wire2(163, 6)    <= sub_wire94(6);
	sub_wire2(163, 7)    <= sub_wire94(7);
	sub_wire2(162, 0)    <= sub_wire95(0);
	sub_wire2(162, 1)    <= sub_wire95(1);
	sub_wire2(162, 2)    <= sub_wire95(2);
	sub_wire2(162, 3)    <= sub_wire95(3);
	sub_wire2(162, 4)    <= sub_wire95(4);
	sub_wire2(162, 5)    <= sub_wire95(5);
	sub_wire2(162, 6)    <= sub_wire95(6);
	sub_wire2(162, 7)    <= sub_wire95(7);
	sub_wire2(161, 0)    <= sub_wire96(0);
	sub_wire2(161, 1)    <= sub_wire96(1);
	sub_wire2(161, 2)    <= sub_wire96(2);
	sub_wire2(161, 3)    <= sub_wire96(3);
	sub_wire2(161, 4)    <= sub_wire96(4);
	sub_wire2(161, 5)    <= sub_wire96(5);
	sub_wire2(161, 6)    <= sub_wire96(6);
	sub_wire2(161, 7)    <= sub_wire96(7);
	sub_wire2(160, 0)    <= sub_wire97(0);
	sub_wire2(160, 1)    <= sub_wire97(1);
	sub_wire2(160, 2)    <= sub_wire97(2);
	sub_wire2(160, 3)    <= sub_wire97(3);
	sub_wire2(160, 4)    <= sub_wire97(4);
	sub_wire2(160, 5)    <= sub_wire97(5);
	sub_wire2(160, 6)    <= sub_wire97(6);
	sub_wire2(160, 7)    <= sub_wire97(7);
	sub_wire2(159, 0)    <= sub_wire98(0);
	sub_wire2(159, 1)    <= sub_wire98(1);
	sub_wire2(159, 2)    <= sub_wire98(2);
	sub_wire2(159, 3)    <= sub_wire98(3);
	sub_wire2(159, 4)    <= sub_wire98(4);
	sub_wire2(159, 5)    <= sub_wire98(5);
	sub_wire2(159, 6)    <= sub_wire98(6);
	sub_wire2(159, 7)    <= sub_wire98(7);
	sub_wire2(158, 0)    <= sub_wire99(0);
	sub_wire2(158, 1)    <= sub_wire99(1);
	sub_wire2(158, 2)    <= sub_wire99(2);
	sub_wire2(158, 3)    <= sub_wire99(3);
	sub_wire2(158, 4)    <= sub_wire99(4);
	sub_wire2(158, 5)    <= sub_wire99(5);
	sub_wire2(158, 6)    <= sub_wire99(6);
	sub_wire2(158, 7)    <= sub_wire99(7);
	sub_wire2(157, 0)    <= sub_wire100(0);
	sub_wire2(157, 1)    <= sub_wire100(1);
	sub_wire2(157, 2)    <= sub_wire100(2);
	sub_wire2(157, 3)    <= sub_wire100(3);
	sub_wire2(157, 4)    <= sub_wire100(4);
	sub_wire2(157, 5)    <= sub_wire100(5);
	sub_wire2(157, 6)    <= sub_wire100(6);
	sub_wire2(157, 7)    <= sub_wire100(7);
	sub_wire2(156, 0)    <= sub_wire101(0);
	sub_wire2(156, 1)    <= sub_wire101(1);
	sub_wire2(156, 2)    <= sub_wire101(2);
	sub_wire2(156, 3)    <= sub_wire101(3);
	sub_wire2(156, 4)    <= sub_wire101(4);
	sub_wire2(156, 5)    <= sub_wire101(5);
	sub_wire2(156, 6)    <= sub_wire101(6);
	sub_wire2(156, 7)    <= sub_wire101(7);
	sub_wire2(155, 0)    <= sub_wire102(0);
	sub_wire2(155, 1)    <= sub_wire102(1);
	sub_wire2(155, 2)    <= sub_wire102(2);
	sub_wire2(155, 3)    <= sub_wire102(3);
	sub_wire2(155, 4)    <= sub_wire102(4);
	sub_wire2(155, 5)    <= sub_wire102(5);
	sub_wire2(155, 6)    <= sub_wire102(6);
	sub_wire2(155, 7)    <= sub_wire102(7);
	sub_wire2(154, 0)    <= sub_wire103(0);
	sub_wire2(154, 1)    <= sub_wire103(1);
	sub_wire2(154, 2)    <= sub_wire103(2);
	sub_wire2(154, 3)    <= sub_wire103(3);
	sub_wire2(154, 4)    <= sub_wire103(4);
	sub_wire2(154, 5)    <= sub_wire103(5);
	sub_wire2(154, 6)    <= sub_wire103(6);
	sub_wire2(154, 7)    <= sub_wire103(7);
	sub_wire2(153, 0)    <= sub_wire104(0);
	sub_wire2(153, 1)    <= sub_wire104(1);
	sub_wire2(153, 2)    <= sub_wire104(2);
	sub_wire2(153, 3)    <= sub_wire104(3);
	sub_wire2(153, 4)    <= sub_wire104(4);
	sub_wire2(153, 5)    <= sub_wire104(5);
	sub_wire2(153, 6)    <= sub_wire104(6);
	sub_wire2(153, 7)    <= sub_wire104(7);
	sub_wire2(152, 0)    <= sub_wire105(0);
	sub_wire2(152, 1)    <= sub_wire105(1);
	sub_wire2(152, 2)    <= sub_wire105(2);
	sub_wire2(152, 3)    <= sub_wire105(3);
	sub_wire2(152, 4)    <= sub_wire105(4);
	sub_wire2(152, 5)    <= sub_wire105(5);
	sub_wire2(152, 6)    <= sub_wire105(6);
	sub_wire2(152, 7)    <= sub_wire105(7);
	sub_wire2(151, 0)    <= sub_wire106(0);
	sub_wire2(151, 1)    <= sub_wire106(1);
	sub_wire2(151, 2)    <= sub_wire106(2);
	sub_wire2(151, 3)    <= sub_wire106(3);
	sub_wire2(151, 4)    <= sub_wire106(4);
	sub_wire2(151, 5)    <= sub_wire106(5);
	sub_wire2(151, 6)    <= sub_wire106(6);
	sub_wire2(151, 7)    <= sub_wire106(7);
	sub_wire2(150, 0)    <= sub_wire107(0);
	sub_wire2(150, 1)    <= sub_wire107(1);
	sub_wire2(150, 2)    <= sub_wire107(2);
	sub_wire2(150, 3)    <= sub_wire107(3);
	sub_wire2(150, 4)    <= sub_wire107(4);
	sub_wire2(150, 5)    <= sub_wire107(5);
	sub_wire2(150, 6)    <= sub_wire107(6);
	sub_wire2(150, 7)    <= sub_wire107(7);
	sub_wire2(149, 0)    <= sub_wire108(0);
	sub_wire2(149, 1)    <= sub_wire108(1);
	sub_wire2(149, 2)    <= sub_wire108(2);
	sub_wire2(149, 3)    <= sub_wire108(3);
	sub_wire2(149, 4)    <= sub_wire108(4);
	sub_wire2(149, 5)    <= sub_wire108(5);
	sub_wire2(149, 6)    <= sub_wire108(6);
	sub_wire2(149, 7)    <= sub_wire108(7);
	sub_wire2(148, 0)    <= sub_wire109(0);
	sub_wire2(148, 1)    <= sub_wire109(1);
	sub_wire2(148, 2)    <= sub_wire109(2);
	sub_wire2(148, 3)    <= sub_wire109(3);
	sub_wire2(148, 4)    <= sub_wire109(4);
	sub_wire2(148, 5)    <= sub_wire109(5);
	sub_wire2(148, 6)    <= sub_wire109(6);
	sub_wire2(148, 7)    <= sub_wire109(7);
	sub_wire2(147, 0)    <= sub_wire110(0);
	sub_wire2(147, 1)    <= sub_wire110(1);
	sub_wire2(147, 2)    <= sub_wire110(2);
	sub_wire2(147, 3)    <= sub_wire110(3);
	sub_wire2(147, 4)    <= sub_wire110(4);
	sub_wire2(147, 5)    <= sub_wire110(5);
	sub_wire2(147, 6)    <= sub_wire110(6);
	sub_wire2(147, 7)    <= sub_wire110(7);
	sub_wire2(146, 0)    <= sub_wire111(0);
	sub_wire2(146, 1)    <= sub_wire111(1);
	sub_wire2(146, 2)    <= sub_wire111(2);
	sub_wire2(146, 3)    <= sub_wire111(3);
	sub_wire2(146, 4)    <= sub_wire111(4);
	sub_wire2(146, 5)    <= sub_wire111(5);
	sub_wire2(146, 6)    <= sub_wire111(6);
	sub_wire2(146, 7)    <= sub_wire111(7);
	sub_wire2(145, 0)    <= sub_wire112(0);
	sub_wire2(145, 1)    <= sub_wire112(1);
	sub_wire2(145, 2)    <= sub_wire112(2);
	sub_wire2(145, 3)    <= sub_wire112(3);
	sub_wire2(145, 4)    <= sub_wire112(4);
	sub_wire2(145, 5)    <= sub_wire112(5);
	sub_wire2(145, 6)    <= sub_wire112(6);
	sub_wire2(145, 7)    <= sub_wire112(7);
	sub_wire2(144, 0)    <= sub_wire113(0);
	sub_wire2(144, 1)    <= sub_wire113(1);
	sub_wire2(144, 2)    <= sub_wire113(2);
	sub_wire2(144, 3)    <= sub_wire113(3);
	sub_wire2(144, 4)    <= sub_wire113(4);
	sub_wire2(144, 5)    <= sub_wire113(5);
	sub_wire2(144, 6)    <= sub_wire113(6);
	sub_wire2(144, 7)    <= sub_wire113(7);
	sub_wire2(143, 0)    <= sub_wire114(0);
	sub_wire2(143, 1)    <= sub_wire114(1);
	sub_wire2(143, 2)    <= sub_wire114(2);
	sub_wire2(143, 3)    <= sub_wire114(3);
	sub_wire2(143, 4)    <= sub_wire114(4);
	sub_wire2(143, 5)    <= sub_wire114(5);
	sub_wire2(143, 6)    <= sub_wire114(6);
	sub_wire2(143, 7)    <= sub_wire114(7);
	sub_wire2(142, 0)    <= sub_wire115(0);
	sub_wire2(142, 1)    <= sub_wire115(1);
	sub_wire2(142, 2)    <= sub_wire115(2);
	sub_wire2(142, 3)    <= sub_wire115(3);
	sub_wire2(142, 4)    <= sub_wire115(4);
	sub_wire2(142, 5)    <= sub_wire115(5);
	sub_wire2(142, 6)    <= sub_wire115(6);
	sub_wire2(142, 7)    <= sub_wire115(7);
	sub_wire2(141, 0)    <= sub_wire116(0);
	sub_wire2(141, 1)    <= sub_wire116(1);
	sub_wire2(141, 2)    <= sub_wire116(2);
	sub_wire2(141, 3)    <= sub_wire116(3);
	sub_wire2(141, 4)    <= sub_wire116(4);
	sub_wire2(141, 5)    <= sub_wire116(5);
	sub_wire2(141, 6)    <= sub_wire116(6);
	sub_wire2(141, 7)    <= sub_wire116(7);
	sub_wire2(140, 0)    <= sub_wire117(0);
	sub_wire2(140, 1)    <= sub_wire117(1);
	sub_wire2(140, 2)    <= sub_wire117(2);
	sub_wire2(140, 3)    <= sub_wire117(3);
	sub_wire2(140, 4)    <= sub_wire117(4);
	sub_wire2(140, 5)    <= sub_wire117(5);
	sub_wire2(140, 6)    <= sub_wire117(6);
	sub_wire2(140, 7)    <= sub_wire117(7);
	sub_wire2(139, 0)    <= sub_wire118(0);
	sub_wire2(139, 1)    <= sub_wire118(1);
	sub_wire2(139, 2)    <= sub_wire118(2);
	sub_wire2(139, 3)    <= sub_wire118(3);
	sub_wire2(139, 4)    <= sub_wire118(4);
	sub_wire2(139, 5)    <= sub_wire118(5);
	sub_wire2(139, 6)    <= sub_wire118(6);
	sub_wire2(139, 7)    <= sub_wire118(7);
	sub_wire2(138, 0)    <= sub_wire119(0);
	sub_wire2(138, 1)    <= sub_wire119(1);
	sub_wire2(138, 2)    <= sub_wire119(2);
	sub_wire2(138, 3)    <= sub_wire119(3);
	sub_wire2(138, 4)    <= sub_wire119(4);
	sub_wire2(138, 5)    <= sub_wire119(5);
	sub_wire2(138, 6)    <= sub_wire119(6);
	sub_wire2(138, 7)    <= sub_wire119(7);
	sub_wire2(137, 0)    <= sub_wire120(0);
	sub_wire2(137, 1)    <= sub_wire120(1);
	sub_wire2(137, 2)    <= sub_wire120(2);
	sub_wire2(137, 3)    <= sub_wire120(3);
	sub_wire2(137, 4)    <= sub_wire120(4);
	sub_wire2(137, 5)    <= sub_wire120(5);
	sub_wire2(137, 6)    <= sub_wire120(6);
	sub_wire2(137, 7)    <= sub_wire120(7);
	sub_wire2(136, 0)    <= sub_wire121(0);
	sub_wire2(136, 1)    <= sub_wire121(1);
	sub_wire2(136, 2)    <= sub_wire121(2);
	sub_wire2(136, 3)    <= sub_wire121(3);
	sub_wire2(136, 4)    <= sub_wire121(4);
	sub_wire2(136, 5)    <= sub_wire121(5);
	sub_wire2(136, 6)    <= sub_wire121(6);
	sub_wire2(136, 7)    <= sub_wire121(7);
	sub_wire2(135, 0)    <= sub_wire122(0);
	sub_wire2(135, 1)    <= sub_wire122(1);
	sub_wire2(135, 2)    <= sub_wire122(2);
	sub_wire2(135, 3)    <= sub_wire122(3);
	sub_wire2(135, 4)    <= sub_wire122(4);
	sub_wire2(135, 5)    <= sub_wire122(5);
	sub_wire2(135, 6)    <= sub_wire122(6);
	sub_wire2(135, 7)    <= sub_wire122(7);
	sub_wire2(134, 0)    <= sub_wire123(0);
	sub_wire2(134, 1)    <= sub_wire123(1);
	sub_wire2(134, 2)    <= sub_wire123(2);
	sub_wire2(134, 3)    <= sub_wire123(3);
	sub_wire2(134, 4)    <= sub_wire123(4);
	sub_wire2(134, 5)    <= sub_wire123(5);
	sub_wire2(134, 6)    <= sub_wire123(6);
	sub_wire2(134, 7)    <= sub_wire123(7);
	sub_wire2(133, 0)    <= sub_wire124(0);
	sub_wire2(133, 1)    <= sub_wire124(1);
	sub_wire2(133, 2)    <= sub_wire124(2);
	sub_wire2(133, 3)    <= sub_wire124(3);
	sub_wire2(133, 4)    <= sub_wire124(4);
	sub_wire2(133, 5)    <= sub_wire124(5);
	sub_wire2(133, 6)    <= sub_wire124(6);
	sub_wire2(133, 7)    <= sub_wire124(7);
	sub_wire2(132, 0)    <= sub_wire125(0);
	sub_wire2(132, 1)    <= sub_wire125(1);
	sub_wire2(132, 2)    <= sub_wire125(2);
	sub_wire2(132, 3)    <= sub_wire125(3);
	sub_wire2(132, 4)    <= sub_wire125(4);
	sub_wire2(132, 5)    <= sub_wire125(5);
	sub_wire2(132, 6)    <= sub_wire125(6);
	sub_wire2(132, 7)    <= sub_wire125(7);
	sub_wire2(131, 0)    <= sub_wire126(0);
	sub_wire2(131, 1)    <= sub_wire126(1);
	sub_wire2(131, 2)    <= sub_wire126(2);
	sub_wire2(131, 3)    <= sub_wire126(3);
	sub_wire2(131, 4)    <= sub_wire126(4);
	sub_wire2(131, 5)    <= sub_wire126(5);
	sub_wire2(131, 6)    <= sub_wire126(6);
	sub_wire2(131, 7)    <= sub_wire126(7);
	sub_wire2(130, 0)    <= sub_wire127(0);
	sub_wire2(130, 1)    <= sub_wire127(1);
	sub_wire2(130, 2)    <= sub_wire127(2);
	sub_wire2(130, 3)    <= sub_wire127(3);
	sub_wire2(130, 4)    <= sub_wire127(4);
	sub_wire2(130, 5)    <= sub_wire127(5);
	sub_wire2(130, 6)    <= sub_wire127(6);
	sub_wire2(130, 7)    <= sub_wire127(7);
	sub_wire2(129, 0)    <= sub_wire128(0);
	sub_wire2(129, 1)    <= sub_wire128(1);
	sub_wire2(129, 2)    <= sub_wire128(2);
	sub_wire2(129, 3)    <= sub_wire128(3);
	sub_wire2(129, 4)    <= sub_wire128(4);
	sub_wire2(129, 5)    <= sub_wire128(5);
	sub_wire2(129, 6)    <= sub_wire128(6);
	sub_wire2(129, 7)    <= sub_wire128(7);
	sub_wire2(128, 0)    <= sub_wire129(0);
	sub_wire2(128, 1)    <= sub_wire129(1);
	sub_wire2(128, 2)    <= sub_wire129(2);
	sub_wire2(128, 3)    <= sub_wire129(3);
	sub_wire2(128, 4)    <= sub_wire129(4);
	sub_wire2(128, 5)    <= sub_wire129(5);
	sub_wire2(128, 6)    <= sub_wire129(6);
	sub_wire2(128, 7)    <= sub_wire129(7);
	sub_wire2(127, 0)    <= sub_wire130(0);
	sub_wire2(127, 1)    <= sub_wire130(1);
	sub_wire2(127, 2)    <= sub_wire130(2);
	sub_wire2(127, 3)    <= sub_wire130(3);
	sub_wire2(127, 4)    <= sub_wire130(4);
	sub_wire2(127, 5)    <= sub_wire130(5);
	sub_wire2(127, 6)    <= sub_wire130(6);
	sub_wire2(127, 7)    <= sub_wire130(7);
	sub_wire2(126, 0)    <= sub_wire131(0);
	sub_wire2(126, 1)    <= sub_wire131(1);
	sub_wire2(126, 2)    <= sub_wire131(2);
	sub_wire2(126, 3)    <= sub_wire131(3);
	sub_wire2(126, 4)    <= sub_wire131(4);
	sub_wire2(126, 5)    <= sub_wire131(5);
	sub_wire2(126, 6)    <= sub_wire131(6);
	sub_wire2(126, 7)    <= sub_wire131(7);
	sub_wire2(125, 0)    <= sub_wire132(0);
	sub_wire2(125, 1)    <= sub_wire132(1);
	sub_wire2(125, 2)    <= sub_wire132(2);
	sub_wire2(125, 3)    <= sub_wire132(3);
	sub_wire2(125, 4)    <= sub_wire132(4);
	sub_wire2(125, 5)    <= sub_wire132(5);
	sub_wire2(125, 6)    <= sub_wire132(6);
	sub_wire2(125, 7)    <= sub_wire132(7);
	sub_wire2(124, 0)    <= sub_wire133(0);
	sub_wire2(124, 1)    <= sub_wire133(1);
	sub_wire2(124, 2)    <= sub_wire133(2);
	sub_wire2(124, 3)    <= sub_wire133(3);
	sub_wire2(124, 4)    <= sub_wire133(4);
	sub_wire2(124, 5)    <= sub_wire133(5);
	sub_wire2(124, 6)    <= sub_wire133(6);
	sub_wire2(124, 7)    <= sub_wire133(7);
	sub_wire2(123, 0)    <= sub_wire134(0);
	sub_wire2(123, 1)    <= sub_wire134(1);
	sub_wire2(123, 2)    <= sub_wire134(2);
	sub_wire2(123, 3)    <= sub_wire134(3);
	sub_wire2(123, 4)    <= sub_wire134(4);
	sub_wire2(123, 5)    <= sub_wire134(5);
	sub_wire2(123, 6)    <= sub_wire134(6);
	sub_wire2(123, 7)    <= sub_wire134(7);
	sub_wire2(122, 0)    <= sub_wire135(0);
	sub_wire2(122, 1)    <= sub_wire135(1);
	sub_wire2(122, 2)    <= sub_wire135(2);
	sub_wire2(122, 3)    <= sub_wire135(3);
	sub_wire2(122, 4)    <= sub_wire135(4);
	sub_wire2(122, 5)    <= sub_wire135(5);
	sub_wire2(122, 6)    <= sub_wire135(6);
	sub_wire2(122, 7)    <= sub_wire135(7);
	sub_wire2(121, 0)    <= sub_wire136(0);
	sub_wire2(121, 1)    <= sub_wire136(1);
	sub_wire2(121, 2)    <= sub_wire136(2);
	sub_wire2(121, 3)    <= sub_wire136(3);
	sub_wire2(121, 4)    <= sub_wire136(4);
	sub_wire2(121, 5)    <= sub_wire136(5);
	sub_wire2(121, 6)    <= sub_wire136(6);
	sub_wire2(121, 7)    <= sub_wire136(7);
	sub_wire2(120, 0)    <= sub_wire137(0);
	sub_wire2(120, 1)    <= sub_wire137(1);
	sub_wire2(120, 2)    <= sub_wire137(2);
	sub_wire2(120, 3)    <= sub_wire137(3);
	sub_wire2(120, 4)    <= sub_wire137(4);
	sub_wire2(120, 5)    <= sub_wire137(5);
	sub_wire2(120, 6)    <= sub_wire137(6);
	sub_wire2(120, 7)    <= sub_wire137(7);
	sub_wire2(119, 0)    <= sub_wire138(0);
	sub_wire2(119, 1)    <= sub_wire138(1);
	sub_wire2(119, 2)    <= sub_wire138(2);
	sub_wire2(119, 3)    <= sub_wire138(3);
	sub_wire2(119, 4)    <= sub_wire138(4);
	sub_wire2(119, 5)    <= sub_wire138(5);
	sub_wire2(119, 6)    <= sub_wire138(6);
	sub_wire2(119, 7)    <= sub_wire138(7);
	sub_wire2(118, 0)    <= sub_wire139(0);
	sub_wire2(118, 1)    <= sub_wire139(1);
	sub_wire2(118, 2)    <= sub_wire139(2);
	sub_wire2(118, 3)    <= sub_wire139(3);
	sub_wire2(118, 4)    <= sub_wire139(4);
	sub_wire2(118, 5)    <= sub_wire139(5);
	sub_wire2(118, 6)    <= sub_wire139(6);
	sub_wire2(118, 7)    <= sub_wire139(7);
	sub_wire2(117, 0)    <= sub_wire140(0);
	sub_wire2(117, 1)    <= sub_wire140(1);
	sub_wire2(117, 2)    <= sub_wire140(2);
	sub_wire2(117, 3)    <= sub_wire140(3);
	sub_wire2(117, 4)    <= sub_wire140(4);
	sub_wire2(117, 5)    <= sub_wire140(5);
	sub_wire2(117, 6)    <= sub_wire140(6);
	sub_wire2(117, 7)    <= sub_wire140(7);
	sub_wire2(116, 0)    <= sub_wire141(0);
	sub_wire2(116, 1)    <= sub_wire141(1);
	sub_wire2(116, 2)    <= sub_wire141(2);
	sub_wire2(116, 3)    <= sub_wire141(3);
	sub_wire2(116, 4)    <= sub_wire141(4);
	sub_wire2(116, 5)    <= sub_wire141(5);
	sub_wire2(116, 6)    <= sub_wire141(6);
	sub_wire2(116, 7)    <= sub_wire141(7);
	sub_wire2(115, 0)    <= sub_wire142(0);
	sub_wire2(115, 1)    <= sub_wire142(1);
	sub_wire2(115, 2)    <= sub_wire142(2);
	sub_wire2(115, 3)    <= sub_wire142(3);
	sub_wire2(115, 4)    <= sub_wire142(4);
	sub_wire2(115, 5)    <= sub_wire142(5);
	sub_wire2(115, 6)    <= sub_wire142(6);
	sub_wire2(115, 7)    <= sub_wire142(7);
	sub_wire2(114, 0)    <= sub_wire143(0);
	sub_wire2(114, 1)    <= sub_wire143(1);
	sub_wire2(114, 2)    <= sub_wire143(2);
	sub_wire2(114, 3)    <= sub_wire143(3);
	sub_wire2(114, 4)    <= sub_wire143(4);
	sub_wire2(114, 5)    <= sub_wire143(5);
	sub_wire2(114, 6)    <= sub_wire143(6);
	sub_wire2(114, 7)    <= sub_wire143(7);
	sub_wire2(113, 0)    <= sub_wire144(0);
	sub_wire2(113, 1)    <= sub_wire144(1);
	sub_wire2(113, 2)    <= sub_wire144(2);
	sub_wire2(113, 3)    <= sub_wire144(3);
	sub_wire2(113, 4)    <= sub_wire144(4);
	sub_wire2(113, 5)    <= sub_wire144(5);
	sub_wire2(113, 6)    <= sub_wire144(6);
	sub_wire2(113, 7)    <= sub_wire144(7);
	sub_wire2(112, 0)    <= sub_wire145(0);
	sub_wire2(112, 1)    <= sub_wire145(1);
	sub_wire2(112, 2)    <= sub_wire145(2);
	sub_wire2(112, 3)    <= sub_wire145(3);
	sub_wire2(112, 4)    <= sub_wire145(4);
	sub_wire2(112, 5)    <= sub_wire145(5);
	sub_wire2(112, 6)    <= sub_wire145(6);
	sub_wire2(112, 7)    <= sub_wire145(7);
	sub_wire2(111, 0)    <= sub_wire146(0);
	sub_wire2(111, 1)    <= sub_wire146(1);
	sub_wire2(111, 2)    <= sub_wire146(2);
	sub_wire2(111, 3)    <= sub_wire146(3);
	sub_wire2(111, 4)    <= sub_wire146(4);
	sub_wire2(111, 5)    <= sub_wire146(5);
	sub_wire2(111, 6)    <= sub_wire146(6);
	sub_wire2(111, 7)    <= sub_wire146(7);
	sub_wire2(110, 0)    <= sub_wire147(0);
	sub_wire2(110, 1)    <= sub_wire147(1);
	sub_wire2(110, 2)    <= sub_wire147(2);
	sub_wire2(110, 3)    <= sub_wire147(3);
	sub_wire2(110, 4)    <= sub_wire147(4);
	sub_wire2(110, 5)    <= sub_wire147(5);
	sub_wire2(110, 6)    <= sub_wire147(6);
	sub_wire2(110, 7)    <= sub_wire147(7);
	sub_wire2(109, 0)    <= sub_wire148(0);
	sub_wire2(109, 1)    <= sub_wire148(1);
	sub_wire2(109, 2)    <= sub_wire148(2);
	sub_wire2(109, 3)    <= sub_wire148(3);
	sub_wire2(109, 4)    <= sub_wire148(4);
	sub_wire2(109, 5)    <= sub_wire148(5);
	sub_wire2(109, 6)    <= sub_wire148(6);
	sub_wire2(109, 7)    <= sub_wire148(7);
	sub_wire2(108, 0)    <= sub_wire149(0);
	sub_wire2(108, 1)    <= sub_wire149(1);
	sub_wire2(108, 2)    <= sub_wire149(2);
	sub_wire2(108, 3)    <= sub_wire149(3);
	sub_wire2(108, 4)    <= sub_wire149(4);
	sub_wire2(108, 5)    <= sub_wire149(5);
	sub_wire2(108, 6)    <= sub_wire149(6);
	sub_wire2(108, 7)    <= sub_wire149(7);
	sub_wire2(107, 0)    <= sub_wire150(0);
	sub_wire2(107, 1)    <= sub_wire150(1);
	sub_wire2(107, 2)    <= sub_wire150(2);
	sub_wire2(107, 3)    <= sub_wire150(3);
	sub_wire2(107, 4)    <= sub_wire150(4);
	sub_wire2(107, 5)    <= sub_wire150(5);
	sub_wire2(107, 6)    <= sub_wire150(6);
	sub_wire2(107, 7)    <= sub_wire150(7);
	sub_wire2(106, 0)    <= sub_wire151(0);
	sub_wire2(106, 1)    <= sub_wire151(1);
	sub_wire2(106, 2)    <= sub_wire151(2);
	sub_wire2(106, 3)    <= sub_wire151(3);
	sub_wire2(106, 4)    <= sub_wire151(4);
	sub_wire2(106, 5)    <= sub_wire151(5);
	sub_wire2(106, 6)    <= sub_wire151(6);
	sub_wire2(106, 7)    <= sub_wire151(7);
	sub_wire2(105, 0)    <= sub_wire152(0);
	sub_wire2(105, 1)    <= sub_wire152(1);
	sub_wire2(105, 2)    <= sub_wire152(2);
	sub_wire2(105, 3)    <= sub_wire152(3);
	sub_wire2(105, 4)    <= sub_wire152(4);
	sub_wire2(105, 5)    <= sub_wire152(5);
	sub_wire2(105, 6)    <= sub_wire152(6);
	sub_wire2(105, 7)    <= sub_wire152(7);
	sub_wire2(104, 0)    <= sub_wire153(0);
	sub_wire2(104, 1)    <= sub_wire153(1);
	sub_wire2(104, 2)    <= sub_wire153(2);
	sub_wire2(104, 3)    <= sub_wire153(3);
	sub_wire2(104, 4)    <= sub_wire153(4);
	sub_wire2(104, 5)    <= sub_wire153(5);
	sub_wire2(104, 6)    <= sub_wire153(6);
	sub_wire2(104, 7)    <= sub_wire153(7);
	sub_wire2(103, 0)    <= sub_wire154(0);
	sub_wire2(103, 1)    <= sub_wire154(1);
	sub_wire2(103, 2)    <= sub_wire154(2);
	sub_wire2(103, 3)    <= sub_wire154(3);
	sub_wire2(103, 4)    <= sub_wire154(4);
	sub_wire2(103, 5)    <= sub_wire154(5);
	sub_wire2(103, 6)    <= sub_wire154(6);
	sub_wire2(103, 7)    <= sub_wire154(7);
	sub_wire2(102, 0)    <= sub_wire155(0);
	sub_wire2(102, 1)    <= sub_wire155(1);
	sub_wire2(102, 2)    <= sub_wire155(2);
	sub_wire2(102, 3)    <= sub_wire155(3);
	sub_wire2(102, 4)    <= sub_wire155(4);
	sub_wire2(102, 5)    <= sub_wire155(5);
	sub_wire2(102, 6)    <= sub_wire155(6);
	sub_wire2(102, 7)    <= sub_wire155(7);
	sub_wire2(101, 0)    <= sub_wire156(0);
	sub_wire2(101, 1)    <= sub_wire156(1);
	sub_wire2(101, 2)    <= sub_wire156(2);
	sub_wire2(101, 3)    <= sub_wire156(3);
	sub_wire2(101, 4)    <= sub_wire156(4);
	sub_wire2(101, 5)    <= sub_wire156(5);
	sub_wire2(101, 6)    <= sub_wire156(6);
	sub_wire2(101, 7)    <= sub_wire156(7);
	sub_wire2(100, 0)    <= sub_wire157(0);
	sub_wire2(100, 1)    <= sub_wire157(1);
	sub_wire2(100, 2)    <= sub_wire157(2);
	sub_wire2(100, 3)    <= sub_wire157(3);
	sub_wire2(100, 4)    <= sub_wire157(4);
	sub_wire2(100, 5)    <= sub_wire157(5);
	sub_wire2(100, 6)    <= sub_wire157(6);
	sub_wire2(100, 7)    <= sub_wire157(7);
	sub_wire2(99, 0)    <= sub_wire158(0);
	sub_wire2(99, 1)    <= sub_wire158(1);
	sub_wire2(99, 2)    <= sub_wire158(2);
	sub_wire2(99, 3)    <= sub_wire158(3);
	sub_wire2(99, 4)    <= sub_wire158(4);
	sub_wire2(99, 5)    <= sub_wire158(5);
	sub_wire2(99, 6)    <= sub_wire158(6);
	sub_wire2(99, 7)    <= sub_wire158(7);
	sub_wire2(98, 0)    <= sub_wire159(0);
	sub_wire2(98, 1)    <= sub_wire159(1);
	sub_wire2(98, 2)    <= sub_wire159(2);
	sub_wire2(98, 3)    <= sub_wire159(3);
	sub_wire2(98, 4)    <= sub_wire159(4);
	sub_wire2(98, 5)    <= sub_wire159(5);
	sub_wire2(98, 6)    <= sub_wire159(6);
	sub_wire2(98, 7)    <= sub_wire159(7);
	sub_wire2(97, 0)    <= sub_wire160(0);
	sub_wire2(97, 1)    <= sub_wire160(1);
	sub_wire2(97, 2)    <= sub_wire160(2);
	sub_wire2(97, 3)    <= sub_wire160(3);
	sub_wire2(97, 4)    <= sub_wire160(4);
	sub_wire2(97, 5)    <= sub_wire160(5);
	sub_wire2(97, 6)    <= sub_wire160(6);
	sub_wire2(97, 7)    <= sub_wire160(7);
	sub_wire2(96, 0)    <= sub_wire161(0);
	sub_wire2(96, 1)    <= sub_wire161(1);
	sub_wire2(96, 2)    <= sub_wire161(2);
	sub_wire2(96, 3)    <= sub_wire161(3);
	sub_wire2(96, 4)    <= sub_wire161(4);
	sub_wire2(96, 5)    <= sub_wire161(5);
	sub_wire2(96, 6)    <= sub_wire161(6);
	sub_wire2(96, 7)    <= sub_wire161(7);
	sub_wire2(95, 0)    <= sub_wire162(0);
	sub_wire2(95, 1)    <= sub_wire162(1);
	sub_wire2(95, 2)    <= sub_wire162(2);
	sub_wire2(95, 3)    <= sub_wire162(3);
	sub_wire2(95, 4)    <= sub_wire162(4);
	sub_wire2(95, 5)    <= sub_wire162(5);
	sub_wire2(95, 6)    <= sub_wire162(6);
	sub_wire2(95, 7)    <= sub_wire162(7);
	sub_wire2(94, 0)    <= sub_wire163(0);
	sub_wire2(94, 1)    <= sub_wire163(1);
	sub_wire2(94, 2)    <= sub_wire163(2);
	sub_wire2(94, 3)    <= sub_wire163(3);
	sub_wire2(94, 4)    <= sub_wire163(4);
	sub_wire2(94, 5)    <= sub_wire163(5);
	sub_wire2(94, 6)    <= sub_wire163(6);
	sub_wire2(94, 7)    <= sub_wire163(7);
	sub_wire2(93, 0)    <= sub_wire164(0);
	sub_wire2(93, 1)    <= sub_wire164(1);
	sub_wire2(93, 2)    <= sub_wire164(2);
	sub_wire2(93, 3)    <= sub_wire164(3);
	sub_wire2(93, 4)    <= sub_wire164(4);
	sub_wire2(93, 5)    <= sub_wire164(5);
	sub_wire2(93, 6)    <= sub_wire164(6);
	sub_wire2(93, 7)    <= sub_wire164(7);
	sub_wire2(92, 0)    <= sub_wire165(0);
	sub_wire2(92, 1)    <= sub_wire165(1);
	sub_wire2(92, 2)    <= sub_wire165(2);
	sub_wire2(92, 3)    <= sub_wire165(3);
	sub_wire2(92, 4)    <= sub_wire165(4);
	sub_wire2(92, 5)    <= sub_wire165(5);
	sub_wire2(92, 6)    <= sub_wire165(6);
	sub_wire2(92, 7)    <= sub_wire165(7);
	sub_wire2(91, 0)    <= sub_wire166(0);
	sub_wire2(91, 1)    <= sub_wire166(1);
	sub_wire2(91, 2)    <= sub_wire166(2);
	sub_wire2(91, 3)    <= sub_wire166(3);
	sub_wire2(91, 4)    <= sub_wire166(4);
	sub_wire2(91, 5)    <= sub_wire166(5);
	sub_wire2(91, 6)    <= sub_wire166(6);
	sub_wire2(91, 7)    <= sub_wire166(7);
	sub_wire2(90, 0)    <= sub_wire167(0);
	sub_wire2(90, 1)    <= sub_wire167(1);
	sub_wire2(90, 2)    <= sub_wire167(2);
	sub_wire2(90, 3)    <= sub_wire167(3);
	sub_wire2(90, 4)    <= sub_wire167(4);
	sub_wire2(90, 5)    <= sub_wire167(5);
	sub_wire2(90, 6)    <= sub_wire167(6);
	sub_wire2(90, 7)    <= sub_wire167(7);
	sub_wire2(89, 0)    <= sub_wire168(0);
	sub_wire2(89, 1)    <= sub_wire168(1);
	sub_wire2(89, 2)    <= sub_wire168(2);
	sub_wire2(89, 3)    <= sub_wire168(3);
	sub_wire2(89, 4)    <= sub_wire168(4);
	sub_wire2(89, 5)    <= sub_wire168(5);
	sub_wire2(89, 6)    <= sub_wire168(6);
	sub_wire2(89, 7)    <= sub_wire168(7);
	sub_wire2(88, 0)    <= sub_wire169(0);
	sub_wire2(88, 1)    <= sub_wire169(1);
	sub_wire2(88, 2)    <= sub_wire169(2);
	sub_wire2(88, 3)    <= sub_wire169(3);
	sub_wire2(88, 4)    <= sub_wire169(4);
	sub_wire2(88, 5)    <= sub_wire169(5);
	sub_wire2(88, 6)    <= sub_wire169(6);
	sub_wire2(88, 7)    <= sub_wire169(7);
	sub_wire2(87, 0)    <= sub_wire170(0);
	sub_wire2(87, 1)    <= sub_wire170(1);
	sub_wire2(87, 2)    <= sub_wire170(2);
	sub_wire2(87, 3)    <= sub_wire170(3);
	sub_wire2(87, 4)    <= sub_wire170(4);
	sub_wire2(87, 5)    <= sub_wire170(5);
	sub_wire2(87, 6)    <= sub_wire170(6);
	sub_wire2(87, 7)    <= sub_wire170(7);
	sub_wire2(86, 0)    <= sub_wire171(0);
	sub_wire2(86, 1)    <= sub_wire171(1);
	sub_wire2(86, 2)    <= sub_wire171(2);
	sub_wire2(86, 3)    <= sub_wire171(3);
	sub_wire2(86, 4)    <= sub_wire171(4);
	sub_wire2(86, 5)    <= sub_wire171(5);
	sub_wire2(86, 6)    <= sub_wire171(6);
	sub_wire2(86, 7)    <= sub_wire171(7);
	sub_wire2(85, 0)    <= sub_wire172(0);
	sub_wire2(85, 1)    <= sub_wire172(1);
	sub_wire2(85, 2)    <= sub_wire172(2);
	sub_wire2(85, 3)    <= sub_wire172(3);
	sub_wire2(85, 4)    <= sub_wire172(4);
	sub_wire2(85, 5)    <= sub_wire172(5);
	sub_wire2(85, 6)    <= sub_wire172(6);
	sub_wire2(85, 7)    <= sub_wire172(7);
	sub_wire2(84, 0)    <= sub_wire173(0);
	sub_wire2(84, 1)    <= sub_wire173(1);
	sub_wire2(84, 2)    <= sub_wire173(2);
	sub_wire2(84, 3)    <= sub_wire173(3);
	sub_wire2(84, 4)    <= sub_wire173(4);
	sub_wire2(84, 5)    <= sub_wire173(5);
	sub_wire2(84, 6)    <= sub_wire173(6);
	sub_wire2(84, 7)    <= sub_wire173(7);
	sub_wire2(83, 0)    <= sub_wire174(0);
	sub_wire2(83, 1)    <= sub_wire174(1);
	sub_wire2(83, 2)    <= sub_wire174(2);
	sub_wire2(83, 3)    <= sub_wire174(3);
	sub_wire2(83, 4)    <= sub_wire174(4);
	sub_wire2(83, 5)    <= sub_wire174(5);
	sub_wire2(83, 6)    <= sub_wire174(6);
	sub_wire2(83, 7)    <= sub_wire174(7);
	sub_wire2(82, 0)    <= sub_wire175(0);
	sub_wire2(82, 1)    <= sub_wire175(1);
	sub_wire2(82, 2)    <= sub_wire175(2);
	sub_wire2(82, 3)    <= sub_wire175(3);
	sub_wire2(82, 4)    <= sub_wire175(4);
	sub_wire2(82, 5)    <= sub_wire175(5);
	sub_wire2(82, 6)    <= sub_wire175(6);
	sub_wire2(82, 7)    <= sub_wire175(7);
	sub_wire2(81, 0)    <= sub_wire176(0);
	sub_wire2(81, 1)    <= sub_wire176(1);
	sub_wire2(81, 2)    <= sub_wire176(2);
	sub_wire2(81, 3)    <= sub_wire176(3);
	sub_wire2(81, 4)    <= sub_wire176(4);
	sub_wire2(81, 5)    <= sub_wire176(5);
	sub_wire2(81, 6)    <= sub_wire176(6);
	sub_wire2(81, 7)    <= sub_wire176(7);
	sub_wire2(80, 0)    <= sub_wire177(0);
	sub_wire2(80, 1)    <= sub_wire177(1);
	sub_wire2(80, 2)    <= sub_wire177(2);
	sub_wire2(80, 3)    <= sub_wire177(3);
	sub_wire2(80, 4)    <= sub_wire177(4);
	sub_wire2(80, 5)    <= sub_wire177(5);
	sub_wire2(80, 6)    <= sub_wire177(6);
	sub_wire2(80, 7)    <= sub_wire177(7);
	sub_wire2(79, 0)    <= sub_wire178(0);
	sub_wire2(79, 1)    <= sub_wire178(1);
	sub_wire2(79, 2)    <= sub_wire178(2);
	sub_wire2(79, 3)    <= sub_wire178(3);
	sub_wire2(79, 4)    <= sub_wire178(4);
	sub_wire2(79, 5)    <= sub_wire178(5);
	sub_wire2(79, 6)    <= sub_wire178(6);
	sub_wire2(79, 7)    <= sub_wire178(7);
	sub_wire2(78, 0)    <= sub_wire179(0);
	sub_wire2(78, 1)    <= sub_wire179(1);
	sub_wire2(78, 2)    <= sub_wire179(2);
	sub_wire2(78, 3)    <= sub_wire179(3);
	sub_wire2(78, 4)    <= sub_wire179(4);
	sub_wire2(78, 5)    <= sub_wire179(5);
	sub_wire2(78, 6)    <= sub_wire179(6);
	sub_wire2(78, 7)    <= sub_wire179(7);
	sub_wire2(77, 0)    <= sub_wire180(0);
	sub_wire2(77, 1)    <= sub_wire180(1);
	sub_wire2(77, 2)    <= sub_wire180(2);
	sub_wire2(77, 3)    <= sub_wire180(3);
	sub_wire2(77, 4)    <= sub_wire180(4);
	sub_wire2(77, 5)    <= sub_wire180(5);
	sub_wire2(77, 6)    <= sub_wire180(6);
	sub_wire2(77, 7)    <= sub_wire180(7);
	sub_wire2(76, 0)    <= sub_wire181(0);
	sub_wire2(76, 1)    <= sub_wire181(1);
	sub_wire2(76, 2)    <= sub_wire181(2);
	sub_wire2(76, 3)    <= sub_wire181(3);
	sub_wire2(76, 4)    <= sub_wire181(4);
	sub_wire2(76, 5)    <= sub_wire181(5);
	sub_wire2(76, 6)    <= sub_wire181(6);
	sub_wire2(76, 7)    <= sub_wire181(7);
	sub_wire2(75, 0)    <= sub_wire182(0);
	sub_wire2(75, 1)    <= sub_wire182(1);
	sub_wire2(75, 2)    <= sub_wire182(2);
	sub_wire2(75, 3)    <= sub_wire182(3);
	sub_wire2(75, 4)    <= sub_wire182(4);
	sub_wire2(75, 5)    <= sub_wire182(5);
	sub_wire2(75, 6)    <= sub_wire182(6);
	sub_wire2(75, 7)    <= sub_wire182(7);
	sub_wire2(74, 0)    <= sub_wire183(0);
	sub_wire2(74, 1)    <= sub_wire183(1);
	sub_wire2(74, 2)    <= sub_wire183(2);
	sub_wire2(74, 3)    <= sub_wire183(3);
	sub_wire2(74, 4)    <= sub_wire183(4);
	sub_wire2(74, 5)    <= sub_wire183(5);
	sub_wire2(74, 6)    <= sub_wire183(6);
	sub_wire2(74, 7)    <= sub_wire183(7);
	sub_wire2(73, 0)    <= sub_wire184(0);
	sub_wire2(73, 1)    <= sub_wire184(1);
	sub_wire2(73, 2)    <= sub_wire184(2);
	sub_wire2(73, 3)    <= sub_wire184(3);
	sub_wire2(73, 4)    <= sub_wire184(4);
	sub_wire2(73, 5)    <= sub_wire184(5);
	sub_wire2(73, 6)    <= sub_wire184(6);
	sub_wire2(73, 7)    <= sub_wire184(7);
	sub_wire2(72, 0)    <= sub_wire185(0);
	sub_wire2(72, 1)    <= sub_wire185(1);
	sub_wire2(72, 2)    <= sub_wire185(2);
	sub_wire2(72, 3)    <= sub_wire185(3);
	sub_wire2(72, 4)    <= sub_wire185(4);
	sub_wire2(72, 5)    <= sub_wire185(5);
	sub_wire2(72, 6)    <= sub_wire185(6);
	sub_wire2(72, 7)    <= sub_wire185(7);
	sub_wire2(71, 0)    <= sub_wire186(0);
	sub_wire2(71, 1)    <= sub_wire186(1);
	sub_wire2(71, 2)    <= sub_wire186(2);
	sub_wire2(71, 3)    <= sub_wire186(3);
	sub_wire2(71, 4)    <= sub_wire186(4);
	sub_wire2(71, 5)    <= sub_wire186(5);
	sub_wire2(71, 6)    <= sub_wire186(6);
	sub_wire2(71, 7)    <= sub_wire186(7);
	sub_wire2(70, 0)    <= sub_wire187(0);
	sub_wire2(70, 1)    <= sub_wire187(1);
	sub_wire2(70, 2)    <= sub_wire187(2);
	sub_wire2(70, 3)    <= sub_wire187(3);
	sub_wire2(70, 4)    <= sub_wire187(4);
	sub_wire2(70, 5)    <= sub_wire187(5);
	sub_wire2(70, 6)    <= sub_wire187(6);
	sub_wire2(70, 7)    <= sub_wire187(7);
	sub_wire2(69, 0)    <= sub_wire188(0);
	sub_wire2(69, 1)    <= sub_wire188(1);
	sub_wire2(69, 2)    <= sub_wire188(2);
	sub_wire2(69, 3)    <= sub_wire188(3);
	sub_wire2(69, 4)    <= sub_wire188(4);
	sub_wire2(69, 5)    <= sub_wire188(5);
	sub_wire2(69, 6)    <= sub_wire188(6);
	sub_wire2(69, 7)    <= sub_wire188(7);
	sub_wire2(68, 0)    <= sub_wire189(0);
	sub_wire2(68, 1)    <= sub_wire189(1);
	sub_wire2(68, 2)    <= sub_wire189(2);
	sub_wire2(68, 3)    <= sub_wire189(3);
	sub_wire2(68, 4)    <= sub_wire189(4);
	sub_wire2(68, 5)    <= sub_wire189(5);
	sub_wire2(68, 6)    <= sub_wire189(6);
	sub_wire2(68, 7)    <= sub_wire189(7);
	sub_wire2(67, 0)    <= sub_wire190(0);
	sub_wire2(67, 1)    <= sub_wire190(1);
	sub_wire2(67, 2)    <= sub_wire190(2);
	sub_wire2(67, 3)    <= sub_wire190(3);
	sub_wire2(67, 4)    <= sub_wire190(4);
	sub_wire2(67, 5)    <= sub_wire190(5);
	sub_wire2(67, 6)    <= sub_wire190(6);
	sub_wire2(67, 7)    <= sub_wire190(7);
	sub_wire2(66, 0)    <= sub_wire191(0);
	sub_wire2(66, 1)    <= sub_wire191(1);
	sub_wire2(66, 2)    <= sub_wire191(2);
	sub_wire2(66, 3)    <= sub_wire191(3);
	sub_wire2(66, 4)    <= sub_wire191(4);
	sub_wire2(66, 5)    <= sub_wire191(5);
	sub_wire2(66, 6)    <= sub_wire191(6);
	sub_wire2(66, 7)    <= sub_wire191(7);
	sub_wire2(65, 0)    <= sub_wire192(0);
	sub_wire2(65, 1)    <= sub_wire192(1);
	sub_wire2(65, 2)    <= sub_wire192(2);
	sub_wire2(65, 3)    <= sub_wire192(3);
	sub_wire2(65, 4)    <= sub_wire192(4);
	sub_wire2(65, 5)    <= sub_wire192(5);
	sub_wire2(65, 6)    <= sub_wire192(6);
	sub_wire2(65, 7)    <= sub_wire192(7);
	sub_wire2(64, 0)    <= sub_wire193(0);
	sub_wire2(64, 1)    <= sub_wire193(1);
	sub_wire2(64, 2)    <= sub_wire193(2);
	sub_wire2(64, 3)    <= sub_wire193(3);
	sub_wire2(64, 4)    <= sub_wire193(4);
	sub_wire2(64, 5)    <= sub_wire193(5);
	sub_wire2(64, 6)    <= sub_wire193(6);
	sub_wire2(64, 7)    <= sub_wire193(7);
	sub_wire2(63, 0)    <= sub_wire194(0);
	sub_wire2(63, 1)    <= sub_wire194(1);
	sub_wire2(63, 2)    <= sub_wire194(2);
	sub_wire2(63, 3)    <= sub_wire194(3);
	sub_wire2(63, 4)    <= sub_wire194(4);
	sub_wire2(63, 5)    <= sub_wire194(5);
	sub_wire2(63, 6)    <= sub_wire194(6);
	sub_wire2(63, 7)    <= sub_wire194(7);
	sub_wire2(62, 0)    <= sub_wire195(0);
	sub_wire2(62, 1)    <= sub_wire195(1);
	sub_wire2(62, 2)    <= sub_wire195(2);
	sub_wire2(62, 3)    <= sub_wire195(3);
	sub_wire2(62, 4)    <= sub_wire195(4);
	sub_wire2(62, 5)    <= sub_wire195(5);
	sub_wire2(62, 6)    <= sub_wire195(6);
	sub_wire2(62, 7)    <= sub_wire195(7);
	sub_wire2(61, 0)    <= sub_wire196(0);
	sub_wire2(61, 1)    <= sub_wire196(1);
	sub_wire2(61, 2)    <= sub_wire196(2);
	sub_wire2(61, 3)    <= sub_wire196(3);
	sub_wire2(61, 4)    <= sub_wire196(4);
	sub_wire2(61, 5)    <= sub_wire196(5);
	sub_wire2(61, 6)    <= sub_wire196(6);
	sub_wire2(61, 7)    <= sub_wire196(7);
	sub_wire2(60, 0)    <= sub_wire197(0);
	sub_wire2(60, 1)    <= sub_wire197(1);
	sub_wire2(60, 2)    <= sub_wire197(2);
	sub_wire2(60, 3)    <= sub_wire197(3);
	sub_wire2(60, 4)    <= sub_wire197(4);
	sub_wire2(60, 5)    <= sub_wire197(5);
	sub_wire2(60, 6)    <= sub_wire197(6);
	sub_wire2(60, 7)    <= sub_wire197(7);
	sub_wire2(59, 0)    <= sub_wire198(0);
	sub_wire2(59, 1)    <= sub_wire198(1);
	sub_wire2(59, 2)    <= sub_wire198(2);
	sub_wire2(59, 3)    <= sub_wire198(3);
	sub_wire2(59, 4)    <= sub_wire198(4);
	sub_wire2(59, 5)    <= sub_wire198(5);
	sub_wire2(59, 6)    <= sub_wire198(6);
	sub_wire2(59, 7)    <= sub_wire198(7);
	sub_wire2(58, 0)    <= sub_wire199(0);
	sub_wire2(58, 1)    <= sub_wire199(1);
	sub_wire2(58, 2)    <= sub_wire199(2);
	sub_wire2(58, 3)    <= sub_wire199(3);
	sub_wire2(58, 4)    <= sub_wire199(4);
	sub_wire2(58, 5)    <= sub_wire199(5);
	sub_wire2(58, 6)    <= sub_wire199(6);
	sub_wire2(58, 7)    <= sub_wire199(7);
	sub_wire2(57, 0)    <= sub_wire200(0);
	sub_wire2(57, 1)    <= sub_wire200(1);
	sub_wire2(57, 2)    <= sub_wire200(2);
	sub_wire2(57, 3)    <= sub_wire200(3);
	sub_wire2(57, 4)    <= sub_wire200(4);
	sub_wire2(57, 5)    <= sub_wire200(5);
	sub_wire2(57, 6)    <= sub_wire200(6);
	sub_wire2(57, 7)    <= sub_wire200(7);
	sub_wire2(56, 0)    <= sub_wire201(0);
	sub_wire2(56, 1)    <= sub_wire201(1);
	sub_wire2(56, 2)    <= sub_wire201(2);
	sub_wire2(56, 3)    <= sub_wire201(3);
	sub_wire2(56, 4)    <= sub_wire201(4);
	sub_wire2(56, 5)    <= sub_wire201(5);
	sub_wire2(56, 6)    <= sub_wire201(6);
	sub_wire2(56, 7)    <= sub_wire201(7);
	sub_wire2(55, 0)    <= sub_wire202(0);
	sub_wire2(55, 1)    <= sub_wire202(1);
	sub_wire2(55, 2)    <= sub_wire202(2);
	sub_wire2(55, 3)    <= sub_wire202(3);
	sub_wire2(55, 4)    <= sub_wire202(4);
	sub_wire2(55, 5)    <= sub_wire202(5);
	sub_wire2(55, 6)    <= sub_wire202(6);
	sub_wire2(55, 7)    <= sub_wire202(7);
	sub_wire2(54, 0)    <= sub_wire203(0);
	sub_wire2(54, 1)    <= sub_wire203(1);
	sub_wire2(54, 2)    <= sub_wire203(2);
	sub_wire2(54, 3)    <= sub_wire203(3);
	sub_wire2(54, 4)    <= sub_wire203(4);
	sub_wire2(54, 5)    <= sub_wire203(5);
	sub_wire2(54, 6)    <= sub_wire203(6);
	sub_wire2(54, 7)    <= sub_wire203(7);
	sub_wire2(53, 0)    <= sub_wire204(0);
	sub_wire2(53, 1)    <= sub_wire204(1);
	sub_wire2(53, 2)    <= sub_wire204(2);
	sub_wire2(53, 3)    <= sub_wire204(3);
	sub_wire2(53, 4)    <= sub_wire204(4);
	sub_wire2(53, 5)    <= sub_wire204(5);
	sub_wire2(53, 6)    <= sub_wire204(6);
	sub_wire2(53, 7)    <= sub_wire204(7);
	sub_wire2(52, 0)    <= sub_wire205(0);
	sub_wire2(52, 1)    <= sub_wire205(1);
	sub_wire2(52, 2)    <= sub_wire205(2);
	sub_wire2(52, 3)    <= sub_wire205(3);
	sub_wire2(52, 4)    <= sub_wire205(4);
	sub_wire2(52, 5)    <= sub_wire205(5);
	sub_wire2(52, 6)    <= sub_wire205(6);
	sub_wire2(52, 7)    <= sub_wire205(7);
	sub_wire2(51, 0)    <= sub_wire206(0);
	sub_wire2(51, 1)    <= sub_wire206(1);
	sub_wire2(51, 2)    <= sub_wire206(2);
	sub_wire2(51, 3)    <= sub_wire206(3);
	sub_wire2(51, 4)    <= sub_wire206(4);
	sub_wire2(51, 5)    <= sub_wire206(5);
	sub_wire2(51, 6)    <= sub_wire206(6);
	sub_wire2(51, 7)    <= sub_wire206(7);
	sub_wire2(50, 0)    <= sub_wire207(0);
	sub_wire2(50, 1)    <= sub_wire207(1);
	sub_wire2(50, 2)    <= sub_wire207(2);
	sub_wire2(50, 3)    <= sub_wire207(3);
	sub_wire2(50, 4)    <= sub_wire207(4);
	sub_wire2(50, 5)    <= sub_wire207(5);
	sub_wire2(50, 6)    <= sub_wire207(6);
	sub_wire2(50, 7)    <= sub_wire207(7);
	sub_wire2(49, 0)    <= sub_wire208(0);
	sub_wire2(49, 1)    <= sub_wire208(1);
	sub_wire2(49, 2)    <= sub_wire208(2);
	sub_wire2(49, 3)    <= sub_wire208(3);
	sub_wire2(49, 4)    <= sub_wire208(4);
	sub_wire2(49, 5)    <= sub_wire208(5);
	sub_wire2(49, 6)    <= sub_wire208(6);
	sub_wire2(49, 7)    <= sub_wire208(7);
	sub_wire2(48, 0)    <= sub_wire209(0);
	sub_wire2(48, 1)    <= sub_wire209(1);
	sub_wire2(48, 2)    <= sub_wire209(2);
	sub_wire2(48, 3)    <= sub_wire209(3);
	sub_wire2(48, 4)    <= sub_wire209(4);
	sub_wire2(48, 5)    <= sub_wire209(5);
	sub_wire2(48, 6)    <= sub_wire209(6);
	sub_wire2(48, 7)    <= sub_wire209(7);
	sub_wire2(47, 0)    <= sub_wire210(0);
	sub_wire2(47, 1)    <= sub_wire210(1);
	sub_wire2(47, 2)    <= sub_wire210(2);
	sub_wire2(47, 3)    <= sub_wire210(3);
	sub_wire2(47, 4)    <= sub_wire210(4);
	sub_wire2(47, 5)    <= sub_wire210(5);
	sub_wire2(47, 6)    <= sub_wire210(6);
	sub_wire2(47, 7)    <= sub_wire210(7);
	sub_wire2(46, 0)    <= sub_wire211(0);
	sub_wire2(46, 1)    <= sub_wire211(1);
	sub_wire2(46, 2)    <= sub_wire211(2);
	sub_wire2(46, 3)    <= sub_wire211(3);
	sub_wire2(46, 4)    <= sub_wire211(4);
	sub_wire2(46, 5)    <= sub_wire211(5);
	sub_wire2(46, 6)    <= sub_wire211(6);
	sub_wire2(46, 7)    <= sub_wire211(7);
	sub_wire2(45, 0)    <= sub_wire212(0);
	sub_wire2(45, 1)    <= sub_wire212(1);
	sub_wire2(45, 2)    <= sub_wire212(2);
	sub_wire2(45, 3)    <= sub_wire212(3);
	sub_wire2(45, 4)    <= sub_wire212(4);
	sub_wire2(45, 5)    <= sub_wire212(5);
	sub_wire2(45, 6)    <= sub_wire212(6);
	sub_wire2(45, 7)    <= sub_wire212(7);
	sub_wire2(44, 0)    <= sub_wire213(0);
	sub_wire2(44, 1)    <= sub_wire213(1);
	sub_wire2(44, 2)    <= sub_wire213(2);
	sub_wire2(44, 3)    <= sub_wire213(3);
	sub_wire2(44, 4)    <= sub_wire213(4);
	sub_wire2(44, 5)    <= sub_wire213(5);
	sub_wire2(44, 6)    <= sub_wire213(6);
	sub_wire2(44, 7)    <= sub_wire213(7);
	sub_wire2(43, 0)    <= sub_wire214(0);
	sub_wire2(43, 1)    <= sub_wire214(1);
	sub_wire2(43, 2)    <= sub_wire214(2);
	sub_wire2(43, 3)    <= sub_wire214(3);
	sub_wire2(43, 4)    <= sub_wire214(4);
	sub_wire2(43, 5)    <= sub_wire214(5);
	sub_wire2(43, 6)    <= sub_wire214(6);
	sub_wire2(43, 7)    <= sub_wire214(7);
	sub_wire2(42, 0)    <= sub_wire215(0);
	sub_wire2(42, 1)    <= sub_wire215(1);
	sub_wire2(42, 2)    <= sub_wire215(2);
	sub_wire2(42, 3)    <= sub_wire215(3);
	sub_wire2(42, 4)    <= sub_wire215(4);
	sub_wire2(42, 5)    <= sub_wire215(5);
	sub_wire2(42, 6)    <= sub_wire215(6);
	sub_wire2(42, 7)    <= sub_wire215(7);
	sub_wire2(41, 0)    <= sub_wire216(0);
	sub_wire2(41, 1)    <= sub_wire216(1);
	sub_wire2(41, 2)    <= sub_wire216(2);
	sub_wire2(41, 3)    <= sub_wire216(3);
	sub_wire2(41, 4)    <= sub_wire216(4);
	sub_wire2(41, 5)    <= sub_wire216(5);
	sub_wire2(41, 6)    <= sub_wire216(6);
	sub_wire2(41, 7)    <= sub_wire216(7);
	sub_wire2(40, 0)    <= sub_wire217(0);
	sub_wire2(40, 1)    <= sub_wire217(1);
	sub_wire2(40, 2)    <= sub_wire217(2);
	sub_wire2(40, 3)    <= sub_wire217(3);
	sub_wire2(40, 4)    <= sub_wire217(4);
	sub_wire2(40, 5)    <= sub_wire217(5);
	sub_wire2(40, 6)    <= sub_wire217(6);
	sub_wire2(40, 7)    <= sub_wire217(7);
	sub_wire2(39, 0)    <= sub_wire218(0);
	sub_wire2(39, 1)    <= sub_wire218(1);
	sub_wire2(39, 2)    <= sub_wire218(2);
	sub_wire2(39, 3)    <= sub_wire218(3);
	sub_wire2(39, 4)    <= sub_wire218(4);
	sub_wire2(39, 5)    <= sub_wire218(5);
	sub_wire2(39, 6)    <= sub_wire218(6);
	sub_wire2(39, 7)    <= sub_wire218(7);
	sub_wire2(38, 0)    <= sub_wire219(0);
	sub_wire2(38, 1)    <= sub_wire219(1);
	sub_wire2(38, 2)    <= sub_wire219(2);
	sub_wire2(38, 3)    <= sub_wire219(3);
	sub_wire2(38, 4)    <= sub_wire219(4);
	sub_wire2(38, 5)    <= sub_wire219(5);
	sub_wire2(38, 6)    <= sub_wire219(6);
	sub_wire2(38, 7)    <= sub_wire219(7);
	sub_wire2(37, 0)    <= sub_wire220(0);
	sub_wire2(37, 1)    <= sub_wire220(1);
	sub_wire2(37, 2)    <= sub_wire220(2);
	sub_wire2(37, 3)    <= sub_wire220(3);
	sub_wire2(37, 4)    <= sub_wire220(4);
	sub_wire2(37, 5)    <= sub_wire220(5);
	sub_wire2(37, 6)    <= sub_wire220(6);
	sub_wire2(37, 7)    <= sub_wire220(7);
	sub_wire2(36, 0)    <= sub_wire221(0);
	sub_wire2(36, 1)    <= sub_wire221(1);
	sub_wire2(36, 2)    <= sub_wire221(2);
	sub_wire2(36, 3)    <= sub_wire221(3);
	sub_wire2(36, 4)    <= sub_wire221(4);
	sub_wire2(36, 5)    <= sub_wire221(5);
	sub_wire2(36, 6)    <= sub_wire221(6);
	sub_wire2(36, 7)    <= sub_wire221(7);
	sub_wire2(35, 0)    <= sub_wire222(0);
	sub_wire2(35, 1)    <= sub_wire222(1);
	sub_wire2(35, 2)    <= sub_wire222(2);
	sub_wire2(35, 3)    <= sub_wire222(3);
	sub_wire2(35, 4)    <= sub_wire222(4);
	sub_wire2(35, 5)    <= sub_wire222(5);
	sub_wire2(35, 6)    <= sub_wire222(6);
	sub_wire2(35, 7)    <= sub_wire222(7);
	sub_wire2(34, 0)    <= sub_wire223(0);
	sub_wire2(34, 1)    <= sub_wire223(1);
	sub_wire2(34, 2)    <= sub_wire223(2);
	sub_wire2(34, 3)    <= sub_wire223(3);
	sub_wire2(34, 4)    <= sub_wire223(4);
	sub_wire2(34, 5)    <= sub_wire223(5);
	sub_wire2(34, 6)    <= sub_wire223(6);
	sub_wire2(34, 7)    <= sub_wire223(7);
	sub_wire2(33, 0)    <= sub_wire224(0);
	sub_wire2(33, 1)    <= sub_wire224(1);
	sub_wire2(33, 2)    <= sub_wire224(2);
	sub_wire2(33, 3)    <= sub_wire224(3);
	sub_wire2(33, 4)    <= sub_wire224(4);
	sub_wire2(33, 5)    <= sub_wire224(5);
	sub_wire2(33, 6)    <= sub_wire224(6);
	sub_wire2(33, 7)    <= sub_wire224(7);
	sub_wire2(32, 0)    <= sub_wire225(0);
	sub_wire2(32, 1)    <= sub_wire225(1);
	sub_wire2(32, 2)    <= sub_wire225(2);
	sub_wire2(32, 3)    <= sub_wire225(3);
	sub_wire2(32, 4)    <= sub_wire225(4);
	sub_wire2(32, 5)    <= sub_wire225(5);
	sub_wire2(32, 6)    <= sub_wire225(6);
	sub_wire2(32, 7)    <= sub_wire225(7);
	sub_wire2(31, 0)    <= sub_wire226(0);
	sub_wire2(31, 1)    <= sub_wire226(1);
	sub_wire2(31, 2)    <= sub_wire226(2);
	sub_wire2(31, 3)    <= sub_wire226(3);
	sub_wire2(31, 4)    <= sub_wire226(4);
	sub_wire2(31, 5)    <= sub_wire226(5);
	sub_wire2(31, 6)    <= sub_wire226(6);
	sub_wire2(31, 7)    <= sub_wire226(7);
	sub_wire2(30, 0)    <= sub_wire227(0);
	sub_wire2(30, 1)    <= sub_wire227(1);
	sub_wire2(30, 2)    <= sub_wire227(2);
	sub_wire2(30, 3)    <= sub_wire227(3);
	sub_wire2(30, 4)    <= sub_wire227(4);
	sub_wire2(30, 5)    <= sub_wire227(5);
	sub_wire2(30, 6)    <= sub_wire227(6);
	sub_wire2(30, 7)    <= sub_wire227(7);
	sub_wire2(29, 0)    <= sub_wire228(0);
	sub_wire2(29, 1)    <= sub_wire228(1);
	sub_wire2(29, 2)    <= sub_wire228(2);
	sub_wire2(29, 3)    <= sub_wire228(3);
	sub_wire2(29, 4)    <= sub_wire228(4);
	sub_wire2(29, 5)    <= sub_wire228(5);
	sub_wire2(29, 6)    <= sub_wire228(6);
	sub_wire2(29, 7)    <= sub_wire228(7);
	sub_wire2(28, 0)    <= sub_wire229(0);
	sub_wire2(28, 1)    <= sub_wire229(1);
	sub_wire2(28, 2)    <= sub_wire229(2);
	sub_wire2(28, 3)    <= sub_wire229(3);
	sub_wire2(28, 4)    <= sub_wire229(4);
	sub_wire2(28, 5)    <= sub_wire229(5);
	sub_wire2(28, 6)    <= sub_wire229(6);
	sub_wire2(28, 7)    <= sub_wire229(7);
	sub_wire2(27, 0)    <= sub_wire230(0);
	sub_wire2(27, 1)    <= sub_wire230(1);
	sub_wire2(27, 2)    <= sub_wire230(2);
	sub_wire2(27, 3)    <= sub_wire230(3);
	sub_wire2(27, 4)    <= sub_wire230(4);
	sub_wire2(27, 5)    <= sub_wire230(5);
	sub_wire2(27, 6)    <= sub_wire230(6);
	sub_wire2(27, 7)    <= sub_wire230(7);
	sub_wire2(26, 0)    <= sub_wire231(0);
	sub_wire2(26, 1)    <= sub_wire231(1);
	sub_wire2(26, 2)    <= sub_wire231(2);
	sub_wire2(26, 3)    <= sub_wire231(3);
	sub_wire2(26, 4)    <= sub_wire231(4);
	sub_wire2(26, 5)    <= sub_wire231(5);
	sub_wire2(26, 6)    <= sub_wire231(6);
	sub_wire2(26, 7)    <= sub_wire231(7);
	sub_wire2(25, 0)    <= sub_wire232(0);
	sub_wire2(25, 1)    <= sub_wire232(1);
	sub_wire2(25, 2)    <= sub_wire232(2);
	sub_wire2(25, 3)    <= sub_wire232(3);
	sub_wire2(25, 4)    <= sub_wire232(4);
	sub_wire2(25, 5)    <= sub_wire232(5);
	sub_wire2(25, 6)    <= sub_wire232(6);
	sub_wire2(25, 7)    <= sub_wire232(7);
	sub_wire2(24, 0)    <= sub_wire233(0);
	sub_wire2(24, 1)    <= sub_wire233(1);
	sub_wire2(24, 2)    <= sub_wire233(2);
	sub_wire2(24, 3)    <= sub_wire233(3);
	sub_wire2(24, 4)    <= sub_wire233(4);
	sub_wire2(24, 5)    <= sub_wire233(5);
	sub_wire2(24, 6)    <= sub_wire233(6);
	sub_wire2(24, 7)    <= sub_wire233(7);
	sub_wire2(23, 0)    <= sub_wire234(0);
	sub_wire2(23, 1)    <= sub_wire234(1);
	sub_wire2(23, 2)    <= sub_wire234(2);
	sub_wire2(23, 3)    <= sub_wire234(3);
	sub_wire2(23, 4)    <= sub_wire234(4);
	sub_wire2(23, 5)    <= sub_wire234(5);
	sub_wire2(23, 6)    <= sub_wire234(6);
	sub_wire2(23, 7)    <= sub_wire234(7);
	sub_wire2(22, 0)    <= sub_wire235(0);
	sub_wire2(22, 1)    <= sub_wire235(1);
	sub_wire2(22, 2)    <= sub_wire235(2);
	sub_wire2(22, 3)    <= sub_wire235(3);
	sub_wire2(22, 4)    <= sub_wire235(4);
	sub_wire2(22, 5)    <= sub_wire235(5);
	sub_wire2(22, 6)    <= sub_wire235(6);
	sub_wire2(22, 7)    <= sub_wire235(7);
	sub_wire2(21, 0)    <= sub_wire236(0);
	sub_wire2(21, 1)    <= sub_wire236(1);
	sub_wire2(21, 2)    <= sub_wire236(2);
	sub_wire2(21, 3)    <= sub_wire236(3);
	sub_wire2(21, 4)    <= sub_wire236(4);
	sub_wire2(21, 5)    <= sub_wire236(5);
	sub_wire2(21, 6)    <= sub_wire236(6);
	sub_wire2(21, 7)    <= sub_wire236(7);
	sub_wire2(20, 0)    <= sub_wire237(0);
	sub_wire2(20, 1)    <= sub_wire237(1);
	sub_wire2(20, 2)    <= sub_wire237(2);
	sub_wire2(20, 3)    <= sub_wire237(3);
	sub_wire2(20, 4)    <= sub_wire237(4);
	sub_wire2(20, 5)    <= sub_wire237(5);
	sub_wire2(20, 6)    <= sub_wire237(6);
	sub_wire2(20, 7)    <= sub_wire237(7);
	sub_wire2(19, 0)    <= sub_wire238(0);
	sub_wire2(19, 1)    <= sub_wire238(1);
	sub_wire2(19, 2)    <= sub_wire238(2);
	sub_wire2(19, 3)    <= sub_wire238(3);
	sub_wire2(19, 4)    <= sub_wire238(4);
	sub_wire2(19, 5)    <= sub_wire238(5);
	sub_wire2(19, 6)    <= sub_wire238(6);
	sub_wire2(19, 7)    <= sub_wire238(7);
	sub_wire2(18, 0)    <= sub_wire239(0);
	sub_wire2(18, 1)    <= sub_wire239(1);
	sub_wire2(18, 2)    <= sub_wire239(2);
	sub_wire2(18, 3)    <= sub_wire239(3);
	sub_wire2(18, 4)    <= sub_wire239(4);
	sub_wire2(18, 5)    <= sub_wire239(5);
	sub_wire2(18, 6)    <= sub_wire239(6);
	sub_wire2(18, 7)    <= sub_wire239(7);
	sub_wire2(17, 0)    <= sub_wire240(0);
	sub_wire2(17, 1)    <= sub_wire240(1);
	sub_wire2(17, 2)    <= sub_wire240(2);
	sub_wire2(17, 3)    <= sub_wire240(3);
	sub_wire2(17, 4)    <= sub_wire240(4);
	sub_wire2(17, 5)    <= sub_wire240(5);
	sub_wire2(17, 6)    <= sub_wire240(6);
	sub_wire2(17, 7)    <= sub_wire240(7);
	sub_wire2(16, 0)    <= sub_wire241(0);
	sub_wire2(16, 1)    <= sub_wire241(1);
	sub_wire2(16, 2)    <= sub_wire241(2);
	sub_wire2(16, 3)    <= sub_wire241(3);
	sub_wire2(16, 4)    <= sub_wire241(4);
	sub_wire2(16, 5)    <= sub_wire241(5);
	sub_wire2(16, 6)    <= sub_wire241(6);
	sub_wire2(16, 7)    <= sub_wire241(7);
	sub_wire2(15, 0)    <= sub_wire242(0);
	sub_wire2(15, 1)    <= sub_wire242(1);
	sub_wire2(15, 2)    <= sub_wire242(2);
	sub_wire2(15, 3)    <= sub_wire242(3);
	sub_wire2(15, 4)    <= sub_wire242(4);
	sub_wire2(15, 5)    <= sub_wire242(5);
	sub_wire2(15, 6)    <= sub_wire242(6);
	sub_wire2(15, 7)    <= sub_wire242(7);
	sub_wire2(14, 0)    <= sub_wire243(0);
	sub_wire2(14, 1)    <= sub_wire243(1);
	sub_wire2(14, 2)    <= sub_wire243(2);
	sub_wire2(14, 3)    <= sub_wire243(3);
	sub_wire2(14, 4)    <= sub_wire243(4);
	sub_wire2(14, 5)    <= sub_wire243(5);
	sub_wire2(14, 6)    <= sub_wire243(6);
	sub_wire2(14, 7)    <= sub_wire243(7);
	sub_wire2(13, 0)    <= sub_wire244(0);
	sub_wire2(13, 1)    <= sub_wire244(1);
	sub_wire2(13, 2)    <= sub_wire244(2);
	sub_wire2(13, 3)    <= sub_wire244(3);
	sub_wire2(13, 4)    <= sub_wire244(4);
	sub_wire2(13, 5)    <= sub_wire244(5);
	sub_wire2(13, 6)    <= sub_wire244(6);
	sub_wire2(13, 7)    <= sub_wire244(7);
	sub_wire2(12, 0)    <= sub_wire245(0);
	sub_wire2(12, 1)    <= sub_wire245(1);
	sub_wire2(12, 2)    <= sub_wire245(2);
	sub_wire2(12, 3)    <= sub_wire245(3);
	sub_wire2(12, 4)    <= sub_wire245(4);
	sub_wire2(12, 5)    <= sub_wire245(5);
	sub_wire2(12, 6)    <= sub_wire245(6);
	sub_wire2(12, 7)    <= sub_wire245(7);
	sub_wire2(11, 0)    <= sub_wire246(0);
	sub_wire2(11, 1)    <= sub_wire246(1);
	sub_wire2(11, 2)    <= sub_wire246(2);
	sub_wire2(11, 3)    <= sub_wire246(3);
	sub_wire2(11, 4)    <= sub_wire246(4);
	sub_wire2(11, 5)    <= sub_wire246(5);
	sub_wire2(11, 6)    <= sub_wire246(6);
	sub_wire2(11, 7)    <= sub_wire246(7);
	sub_wire2(10, 0)    <= sub_wire247(0);
	sub_wire2(10, 1)    <= sub_wire247(1);
	sub_wire2(10, 2)    <= sub_wire247(2);
	sub_wire2(10, 3)    <= sub_wire247(3);
	sub_wire2(10, 4)    <= sub_wire247(4);
	sub_wire2(10, 5)    <= sub_wire247(5);
	sub_wire2(10, 6)    <= sub_wire247(6);
	sub_wire2(10, 7)    <= sub_wire247(7);
	sub_wire2(9, 0)    <= sub_wire248(0);
	sub_wire2(9, 1)    <= sub_wire248(1);
	sub_wire2(9, 2)    <= sub_wire248(2);
	sub_wire2(9, 3)    <= sub_wire248(3);
	sub_wire2(9, 4)    <= sub_wire248(4);
	sub_wire2(9, 5)    <= sub_wire248(5);
	sub_wire2(9, 6)    <= sub_wire248(6);
	sub_wire2(9, 7)    <= sub_wire248(7);
	sub_wire2(8, 0)    <= sub_wire249(0);
	sub_wire2(8, 1)    <= sub_wire249(1);
	sub_wire2(8, 2)    <= sub_wire249(2);
	sub_wire2(8, 3)    <= sub_wire249(3);
	sub_wire2(8, 4)    <= sub_wire249(4);
	sub_wire2(8, 5)    <= sub_wire249(5);
	sub_wire2(8, 6)    <= sub_wire249(6);
	sub_wire2(8, 7)    <= sub_wire249(7);
	sub_wire2(7, 0)    <= sub_wire250(0);
	sub_wire2(7, 1)    <= sub_wire250(1);
	sub_wire2(7, 2)    <= sub_wire250(2);
	sub_wire2(7, 3)    <= sub_wire250(3);
	sub_wire2(7, 4)    <= sub_wire250(4);
	sub_wire2(7, 5)    <= sub_wire250(5);
	sub_wire2(7, 6)    <= sub_wire250(6);
	sub_wire2(7, 7)    <= sub_wire250(7);
	sub_wire2(6, 0)    <= sub_wire251(0);
	sub_wire2(6, 1)    <= sub_wire251(1);
	sub_wire2(6, 2)    <= sub_wire251(2);
	sub_wire2(6, 3)    <= sub_wire251(3);
	sub_wire2(6, 4)    <= sub_wire251(4);
	sub_wire2(6, 5)    <= sub_wire251(5);
	sub_wire2(6, 6)    <= sub_wire251(6);
	sub_wire2(6, 7)    <= sub_wire251(7);
	sub_wire2(5, 0)    <= sub_wire252(0);
	sub_wire2(5, 1)    <= sub_wire252(1);
	sub_wire2(5, 2)    <= sub_wire252(2);
	sub_wire2(5, 3)    <= sub_wire252(3);
	sub_wire2(5, 4)    <= sub_wire252(4);
	sub_wire2(5, 5)    <= sub_wire252(5);
	sub_wire2(5, 6)    <= sub_wire252(6);
	sub_wire2(5, 7)    <= sub_wire252(7);
	sub_wire2(4, 0)    <= sub_wire253(0);
	sub_wire2(4, 1)    <= sub_wire253(1);
	sub_wire2(4, 2)    <= sub_wire253(2);
	sub_wire2(4, 3)    <= sub_wire253(3);
	sub_wire2(4, 4)    <= sub_wire253(4);
	sub_wire2(4, 5)    <= sub_wire253(5);
	sub_wire2(4, 6)    <= sub_wire253(6);
	sub_wire2(4, 7)    <= sub_wire253(7);
	sub_wire2(3, 0)    <= sub_wire254(0);
	sub_wire2(3, 1)    <= sub_wire254(1);
	sub_wire2(3, 2)    <= sub_wire254(2);
	sub_wire2(3, 3)    <= sub_wire254(3);
	sub_wire2(3, 4)    <= sub_wire254(4);
	sub_wire2(3, 5)    <= sub_wire254(5);
	sub_wire2(3, 6)    <= sub_wire254(6);
	sub_wire2(3, 7)    <= sub_wire254(7);
	sub_wire2(2, 0)    <= sub_wire255(0);
	sub_wire2(2, 1)    <= sub_wire255(1);
	sub_wire2(2, 2)    <= sub_wire255(2);
	sub_wire2(2, 3)    <= sub_wire255(3);
	sub_wire2(2, 4)    <= sub_wire255(4);
	sub_wire2(2, 5)    <= sub_wire255(5);
	sub_wire2(2, 6)    <= sub_wire255(6);
	sub_wire2(2, 7)    <= sub_wire255(7);
	sub_wire2(1, 0)    <= sub_wire256(0);
	sub_wire2(1, 1)    <= sub_wire256(1);
	sub_wire2(1, 2)    <= sub_wire256(2);
	sub_wire2(1, 3)    <= sub_wire256(3);
	sub_wire2(1, 4)    <= sub_wire256(4);
	sub_wire2(1, 5)    <= sub_wire256(5);
	sub_wire2(1, 6)    <= sub_wire256(6);
	sub_wire2(1, 7)    <= sub_wire256(7);
	sub_wire2(0, 0)    <= sub_wire257(0);
	sub_wire2(0, 1)    <= sub_wire257(1);
	sub_wire2(0, 2)    <= sub_wire257(2);
	sub_wire2(0, 3)    <= sub_wire257(3);
	sub_wire2(0, 4)    <= sub_wire257(4);
	sub_wire2(0, 5)    <= sub_wire257(5);
	sub_wire2(0, 6)    <= sub_wire257(6);
	sub_wire2(0, 7)    <= sub_wire257(7);

	lpm_mux_component : lpm_mux
	GENERIC MAP (
		lpm_size => 256,
		lpm_type => "LPM_MUX",
		lpm_width => 8,
		lpm_widths => 8
	)
	PORT MAP (
		sel => sel,
		data => sub_wire2,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "256"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "8"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "8"
-- Retrieval info: USED_PORT: data0x 0 0 8 0 INPUT NODEFVAL data0x[7..0]
-- Retrieval info: USED_PORT: data100x 0 0 8 0 INPUT NODEFVAL data100x[7..0]
-- Retrieval info: USED_PORT: data101x 0 0 8 0 INPUT NODEFVAL data101x[7..0]
-- Retrieval info: USED_PORT: data102x 0 0 8 0 INPUT NODEFVAL data102x[7..0]
-- Retrieval info: USED_PORT: data103x 0 0 8 0 INPUT NODEFVAL data103x[7..0]
-- Retrieval info: USED_PORT: data104x 0 0 8 0 INPUT NODEFVAL data104x[7..0]
-- Retrieval info: USED_PORT: data105x 0 0 8 0 INPUT NODEFVAL data105x[7..0]
-- Retrieval info: USED_PORT: data106x 0 0 8 0 INPUT NODEFVAL data106x[7..0]
-- Retrieval info: USED_PORT: data107x 0 0 8 0 INPUT NODEFVAL data107x[7..0]
-- Retrieval info: USED_PORT: data108x 0 0 8 0 INPUT NODEFVAL data108x[7..0]
-- Retrieval info: USED_PORT: data109x 0 0 8 0 INPUT NODEFVAL data109x[7..0]
-- Retrieval info: USED_PORT: data10x 0 0 8 0 INPUT NODEFVAL data10x[7..0]
-- Retrieval info: USED_PORT: data110x 0 0 8 0 INPUT NODEFVAL data110x[7..0]
-- Retrieval info: USED_PORT: data111x 0 0 8 0 INPUT NODEFVAL data111x[7..0]
-- Retrieval info: USED_PORT: data112x 0 0 8 0 INPUT NODEFVAL data112x[7..0]
-- Retrieval info: USED_PORT: data113x 0 0 8 0 INPUT NODEFVAL data113x[7..0]
-- Retrieval info: USED_PORT: data114x 0 0 8 0 INPUT NODEFVAL data114x[7..0]
-- Retrieval info: USED_PORT: data115x 0 0 8 0 INPUT NODEFVAL data115x[7..0]
-- Retrieval info: USED_PORT: data116x 0 0 8 0 INPUT NODEFVAL data116x[7..0]
-- Retrieval info: USED_PORT: data117x 0 0 8 0 INPUT NODEFVAL data117x[7..0]
-- Retrieval info: USED_PORT: data118x 0 0 8 0 INPUT NODEFVAL data118x[7..0]
-- Retrieval info: USED_PORT: data119x 0 0 8 0 INPUT NODEFVAL data119x[7..0]
-- Retrieval info: USED_PORT: data11x 0 0 8 0 INPUT NODEFVAL data11x[7..0]
-- Retrieval info: USED_PORT: data120x 0 0 8 0 INPUT NODEFVAL data120x[7..0]
-- Retrieval info: USED_PORT: data121x 0 0 8 0 INPUT NODEFVAL data121x[7..0]
-- Retrieval info: USED_PORT: data122x 0 0 8 0 INPUT NODEFVAL data122x[7..0]
-- Retrieval info: USED_PORT: data123x 0 0 8 0 INPUT NODEFVAL data123x[7..0]
-- Retrieval info: USED_PORT: data124x 0 0 8 0 INPUT NODEFVAL data124x[7..0]
-- Retrieval info: USED_PORT: data125x 0 0 8 0 INPUT NODEFVAL data125x[7..0]
-- Retrieval info: USED_PORT: data126x 0 0 8 0 INPUT NODEFVAL data126x[7..0]
-- Retrieval info: USED_PORT: data127x 0 0 8 0 INPUT NODEFVAL data127x[7..0]
-- Retrieval info: USED_PORT: data128x 0 0 8 0 INPUT NODEFVAL data128x[7..0]
-- Retrieval info: USED_PORT: data129x 0 0 8 0 INPUT NODEFVAL data129x[7..0]
-- Retrieval info: USED_PORT: data12x 0 0 8 0 INPUT NODEFVAL data12x[7..0]
-- Retrieval info: USED_PORT: data130x 0 0 8 0 INPUT NODEFVAL data130x[7..0]
-- Retrieval info: USED_PORT: data131x 0 0 8 0 INPUT NODEFVAL data131x[7..0]
-- Retrieval info: USED_PORT: data132x 0 0 8 0 INPUT NODEFVAL data132x[7..0]
-- Retrieval info: USED_PORT: data133x 0 0 8 0 INPUT NODEFVAL data133x[7..0]
-- Retrieval info: USED_PORT: data134x 0 0 8 0 INPUT NODEFVAL data134x[7..0]
-- Retrieval info: USED_PORT: data135x 0 0 8 0 INPUT NODEFVAL data135x[7..0]
-- Retrieval info: USED_PORT: data136x 0 0 8 0 INPUT NODEFVAL data136x[7..0]
-- Retrieval info: USED_PORT: data137x 0 0 8 0 INPUT NODEFVAL data137x[7..0]
-- Retrieval info: USED_PORT: data138x 0 0 8 0 INPUT NODEFVAL data138x[7..0]
-- Retrieval info: USED_PORT: data139x 0 0 8 0 INPUT NODEFVAL data139x[7..0]
-- Retrieval info: USED_PORT: data13x 0 0 8 0 INPUT NODEFVAL data13x[7..0]
-- Retrieval info: USED_PORT: data140x 0 0 8 0 INPUT NODEFVAL data140x[7..0]
-- Retrieval info: USED_PORT: data141x 0 0 8 0 INPUT NODEFVAL data141x[7..0]
-- Retrieval info: USED_PORT: data142x 0 0 8 0 INPUT NODEFVAL data142x[7..0]
-- Retrieval info: USED_PORT: data143x 0 0 8 0 INPUT NODEFVAL data143x[7..0]
-- Retrieval info: USED_PORT: data144x 0 0 8 0 INPUT NODEFVAL data144x[7..0]
-- Retrieval info: USED_PORT: data145x 0 0 8 0 INPUT NODEFVAL data145x[7..0]
-- Retrieval info: USED_PORT: data146x 0 0 8 0 INPUT NODEFVAL data146x[7..0]
-- Retrieval info: USED_PORT: data147x 0 0 8 0 INPUT NODEFVAL data147x[7..0]
-- Retrieval info: USED_PORT: data148x 0 0 8 0 INPUT NODEFVAL data148x[7..0]
-- Retrieval info: USED_PORT: data149x 0 0 8 0 INPUT NODEFVAL data149x[7..0]
-- Retrieval info: USED_PORT: data14x 0 0 8 0 INPUT NODEFVAL data14x[7..0]
-- Retrieval info: USED_PORT: data150x 0 0 8 0 INPUT NODEFVAL data150x[7..0]
-- Retrieval info: USED_PORT: data151x 0 0 8 0 INPUT NODEFVAL data151x[7..0]
-- Retrieval info: USED_PORT: data152x 0 0 8 0 INPUT NODEFVAL data152x[7..0]
-- Retrieval info: USED_PORT: data153x 0 0 8 0 INPUT NODEFVAL data153x[7..0]
-- Retrieval info: USED_PORT: data154x 0 0 8 0 INPUT NODEFVAL data154x[7..0]
-- Retrieval info: USED_PORT: data155x 0 0 8 0 INPUT NODEFVAL data155x[7..0]
-- Retrieval info: USED_PORT: data156x 0 0 8 0 INPUT NODEFVAL data156x[7..0]
-- Retrieval info: USED_PORT: data157x 0 0 8 0 INPUT NODEFVAL data157x[7..0]
-- Retrieval info: USED_PORT: data158x 0 0 8 0 INPUT NODEFVAL data158x[7..0]
-- Retrieval info: USED_PORT: data159x 0 0 8 0 INPUT NODEFVAL data159x[7..0]
-- Retrieval info: USED_PORT: data15x 0 0 8 0 INPUT NODEFVAL data15x[7..0]
-- Retrieval info: USED_PORT: data160x 0 0 8 0 INPUT NODEFVAL data160x[7..0]
-- Retrieval info: USED_PORT: data161x 0 0 8 0 INPUT NODEFVAL data161x[7..0]
-- Retrieval info: USED_PORT: data162x 0 0 8 0 INPUT NODEFVAL data162x[7..0]
-- Retrieval info: USED_PORT: data163x 0 0 8 0 INPUT NODEFVAL data163x[7..0]
-- Retrieval info: USED_PORT: data164x 0 0 8 0 INPUT NODEFVAL data164x[7..0]
-- Retrieval info: USED_PORT: data165x 0 0 8 0 INPUT NODEFVAL data165x[7..0]
-- Retrieval info: USED_PORT: data166x 0 0 8 0 INPUT NODEFVAL data166x[7..0]
-- Retrieval info: USED_PORT: data167x 0 0 8 0 INPUT NODEFVAL data167x[7..0]
-- Retrieval info: USED_PORT: data168x 0 0 8 0 INPUT NODEFVAL data168x[7..0]
-- Retrieval info: USED_PORT: data169x 0 0 8 0 INPUT NODEFVAL data169x[7..0]
-- Retrieval info: USED_PORT: data16x 0 0 8 0 INPUT NODEFVAL data16x[7..0]
-- Retrieval info: USED_PORT: data170x 0 0 8 0 INPUT NODEFVAL data170x[7..0]
-- Retrieval info: USED_PORT: data171x 0 0 8 0 INPUT NODEFVAL data171x[7..0]
-- Retrieval info: USED_PORT: data172x 0 0 8 0 INPUT NODEFVAL data172x[7..0]
-- Retrieval info: USED_PORT: data173x 0 0 8 0 INPUT NODEFVAL data173x[7..0]
-- Retrieval info: USED_PORT: data174x 0 0 8 0 INPUT NODEFVAL data174x[7..0]
-- Retrieval info: USED_PORT: data175x 0 0 8 0 INPUT NODEFVAL data175x[7..0]
-- Retrieval info: USED_PORT: data176x 0 0 8 0 INPUT NODEFVAL data176x[7..0]
-- Retrieval info: USED_PORT: data177x 0 0 8 0 INPUT NODEFVAL data177x[7..0]
-- Retrieval info: USED_PORT: data178x 0 0 8 0 INPUT NODEFVAL data178x[7..0]
-- Retrieval info: USED_PORT: data179x 0 0 8 0 INPUT NODEFVAL data179x[7..0]
-- Retrieval info: USED_PORT: data17x 0 0 8 0 INPUT NODEFVAL data17x[7..0]
-- Retrieval info: USED_PORT: data180x 0 0 8 0 INPUT NODEFVAL data180x[7..0]
-- Retrieval info: USED_PORT: data181x 0 0 8 0 INPUT NODEFVAL data181x[7..0]
-- Retrieval info: USED_PORT: data182x 0 0 8 0 INPUT NODEFVAL data182x[7..0]
-- Retrieval info: USED_PORT: data183x 0 0 8 0 INPUT NODEFVAL data183x[7..0]
-- Retrieval info: USED_PORT: data184x 0 0 8 0 INPUT NODEFVAL data184x[7..0]
-- Retrieval info: USED_PORT: data185x 0 0 8 0 INPUT NODEFVAL data185x[7..0]
-- Retrieval info: USED_PORT: data186x 0 0 8 0 INPUT NODEFVAL data186x[7..0]
-- Retrieval info: USED_PORT: data187x 0 0 8 0 INPUT NODEFVAL data187x[7..0]
-- Retrieval info: USED_PORT: data188x 0 0 8 0 INPUT NODEFVAL data188x[7..0]
-- Retrieval info: USED_PORT: data189x 0 0 8 0 INPUT NODEFVAL data189x[7..0]
-- Retrieval info: USED_PORT: data18x 0 0 8 0 INPUT NODEFVAL data18x[7..0]
-- Retrieval info: USED_PORT: data190x 0 0 8 0 INPUT NODEFVAL data190x[7..0]
-- Retrieval info: USED_PORT: data191x 0 0 8 0 INPUT NODEFVAL data191x[7..0]
-- Retrieval info: USED_PORT: data192x 0 0 8 0 INPUT NODEFVAL data192x[7..0]
-- Retrieval info: USED_PORT: data193x 0 0 8 0 INPUT NODEFVAL data193x[7..0]
-- Retrieval info: USED_PORT: data194x 0 0 8 0 INPUT NODEFVAL data194x[7..0]
-- Retrieval info: USED_PORT: data195x 0 0 8 0 INPUT NODEFVAL data195x[7..0]
-- Retrieval info: USED_PORT: data196x 0 0 8 0 INPUT NODEFVAL data196x[7..0]
-- Retrieval info: USED_PORT: data197x 0 0 8 0 INPUT NODEFVAL data197x[7..0]
-- Retrieval info: USED_PORT: data198x 0 0 8 0 INPUT NODEFVAL data198x[7..0]
-- Retrieval info: USED_PORT: data199x 0 0 8 0 INPUT NODEFVAL data199x[7..0]
-- Retrieval info: USED_PORT: data19x 0 0 8 0 INPUT NODEFVAL data19x[7..0]
-- Retrieval info: USED_PORT: data1x 0 0 8 0 INPUT NODEFVAL data1x[7..0]
-- Retrieval info: USED_PORT: data200x 0 0 8 0 INPUT NODEFVAL data200x[7..0]
-- Retrieval info: USED_PORT: data201x 0 0 8 0 INPUT NODEFVAL data201x[7..0]
-- Retrieval info: USED_PORT: data202x 0 0 8 0 INPUT NODEFVAL data202x[7..0]
-- Retrieval info: USED_PORT: data203x 0 0 8 0 INPUT NODEFVAL data203x[7..0]
-- Retrieval info: USED_PORT: data204x 0 0 8 0 INPUT NODEFVAL data204x[7..0]
-- Retrieval info: USED_PORT: data205x 0 0 8 0 INPUT NODEFVAL data205x[7..0]
-- Retrieval info: USED_PORT: data206x 0 0 8 0 INPUT NODEFVAL data206x[7..0]
-- Retrieval info: USED_PORT: data207x 0 0 8 0 INPUT NODEFVAL data207x[7..0]
-- Retrieval info: USED_PORT: data208x 0 0 8 0 INPUT NODEFVAL data208x[7..0]
-- Retrieval info: USED_PORT: data209x 0 0 8 0 INPUT NODEFVAL data209x[7..0]
-- Retrieval info: USED_PORT: data20x 0 0 8 0 INPUT NODEFVAL data20x[7..0]
-- Retrieval info: USED_PORT: data210x 0 0 8 0 INPUT NODEFVAL data210x[7..0]
-- Retrieval info: USED_PORT: data211x 0 0 8 0 INPUT NODEFVAL data211x[7..0]
-- Retrieval info: USED_PORT: data212x 0 0 8 0 INPUT NODEFVAL data212x[7..0]
-- Retrieval info: USED_PORT: data213x 0 0 8 0 INPUT NODEFVAL data213x[7..0]
-- Retrieval info: USED_PORT: data214x 0 0 8 0 INPUT NODEFVAL data214x[7..0]
-- Retrieval info: USED_PORT: data215x 0 0 8 0 INPUT NODEFVAL data215x[7..0]
-- Retrieval info: USED_PORT: data216x 0 0 8 0 INPUT NODEFVAL data216x[7..0]
-- Retrieval info: USED_PORT: data217x 0 0 8 0 INPUT NODEFVAL data217x[7..0]
-- Retrieval info: USED_PORT: data218x 0 0 8 0 INPUT NODEFVAL data218x[7..0]
-- Retrieval info: USED_PORT: data219x 0 0 8 0 INPUT NODEFVAL data219x[7..0]
-- Retrieval info: USED_PORT: data21x 0 0 8 0 INPUT NODEFVAL data21x[7..0]
-- Retrieval info: USED_PORT: data220x 0 0 8 0 INPUT NODEFVAL data220x[7..0]
-- Retrieval info: USED_PORT: data221x 0 0 8 0 INPUT NODEFVAL data221x[7..0]
-- Retrieval info: USED_PORT: data222x 0 0 8 0 INPUT NODEFVAL data222x[7..0]
-- Retrieval info: USED_PORT: data223x 0 0 8 0 INPUT NODEFVAL data223x[7..0]
-- Retrieval info: USED_PORT: data224x 0 0 8 0 INPUT NODEFVAL data224x[7..0]
-- Retrieval info: USED_PORT: data225x 0 0 8 0 INPUT NODEFVAL data225x[7..0]
-- Retrieval info: USED_PORT: data226x 0 0 8 0 INPUT NODEFVAL data226x[7..0]
-- Retrieval info: USED_PORT: data227x 0 0 8 0 INPUT NODEFVAL data227x[7..0]
-- Retrieval info: USED_PORT: data228x 0 0 8 0 INPUT NODEFVAL data228x[7..0]
-- Retrieval info: USED_PORT: data229x 0 0 8 0 INPUT NODEFVAL data229x[7..0]
-- Retrieval info: USED_PORT: data22x 0 0 8 0 INPUT NODEFVAL data22x[7..0]
-- Retrieval info: USED_PORT: data230x 0 0 8 0 INPUT NODEFVAL data230x[7..0]
-- Retrieval info: USED_PORT: data231x 0 0 8 0 INPUT NODEFVAL data231x[7..0]
-- Retrieval info: USED_PORT: data232x 0 0 8 0 INPUT NODEFVAL data232x[7..0]
-- Retrieval info: USED_PORT: data233x 0 0 8 0 INPUT NODEFVAL data233x[7..0]
-- Retrieval info: USED_PORT: data234x 0 0 8 0 INPUT NODEFVAL data234x[7..0]
-- Retrieval info: USED_PORT: data235x 0 0 8 0 INPUT NODEFVAL data235x[7..0]
-- Retrieval info: USED_PORT: data236x 0 0 8 0 INPUT NODEFVAL data236x[7..0]
-- Retrieval info: USED_PORT: data237x 0 0 8 0 INPUT NODEFVAL data237x[7..0]
-- Retrieval info: USED_PORT: data238x 0 0 8 0 INPUT NODEFVAL data238x[7..0]
-- Retrieval info: USED_PORT: data239x 0 0 8 0 INPUT NODEFVAL data239x[7..0]
-- Retrieval info: USED_PORT: data23x 0 0 8 0 INPUT NODEFVAL data23x[7..0]
-- Retrieval info: USED_PORT: data240x 0 0 8 0 INPUT NODEFVAL data240x[7..0]
-- Retrieval info: USED_PORT: data241x 0 0 8 0 INPUT NODEFVAL data241x[7..0]
-- Retrieval info: USED_PORT: data242x 0 0 8 0 INPUT NODEFVAL data242x[7..0]
-- Retrieval info: USED_PORT: data243x 0 0 8 0 INPUT NODEFVAL data243x[7..0]
-- Retrieval info: USED_PORT: data244x 0 0 8 0 INPUT NODEFVAL data244x[7..0]
-- Retrieval info: USED_PORT: data245x 0 0 8 0 INPUT NODEFVAL data245x[7..0]
-- Retrieval info: USED_PORT: data246x 0 0 8 0 INPUT NODEFVAL data246x[7..0]
-- Retrieval info: USED_PORT: data247x 0 0 8 0 INPUT NODEFVAL data247x[7..0]
-- Retrieval info: USED_PORT: data248x 0 0 8 0 INPUT NODEFVAL data248x[7..0]
-- Retrieval info: USED_PORT: data249x 0 0 8 0 INPUT NODEFVAL data249x[7..0]
-- Retrieval info: USED_PORT: data24x 0 0 8 0 INPUT NODEFVAL data24x[7..0]
-- Retrieval info: USED_PORT: data250x 0 0 8 0 INPUT NODEFVAL data250x[7..0]
-- Retrieval info: USED_PORT: data251x 0 0 8 0 INPUT NODEFVAL data251x[7..0]
-- Retrieval info: USED_PORT: data252x 0 0 8 0 INPUT NODEFVAL data252x[7..0]
-- Retrieval info: USED_PORT: data253x 0 0 8 0 INPUT NODEFVAL data253x[7..0]
-- Retrieval info: USED_PORT: data254x 0 0 8 0 INPUT NODEFVAL data254x[7..0]
-- Retrieval info: USED_PORT: data255x 0 0 8 0 INPUT NODEFVAL data255x[7..0]
-- Retrieval info: USED_PORT: data25x 0 0 8 0 INPUT NODEFVAL data25x[7..0]
-- Retrieval info: USED_PORT: data26x 0 0 8 0 INPUT NODEFVAL data26x[7..0]
-- Retrieval info: USED_PORT: data27x 0 0 8 0 INPUT NODEFVAL data27x[7..0]
-- Retrieval info: USED_PORT: data28x 0 0 8 0 INPUT NODEFVAL data28x[7..0]
-- Retrieval info: USED_PORT: data29x 0 0 8 0 INPUT NODEFVAL data29x[7..0]
-- Retrieval info: USED_PORT: data2x 0 0 8 0 INPUT NODEFVAL data2x[7..0]
-- Retrieval info: USED_PORT: data30x 0 0 8 0 INPUT NODEFVAL data30x[7..0]
-- Retrieval info: USED_PORT: data31x 0 0 8 0 INPUT NODEFVAL data31x[7..0]
-- Retrieval info: USED_PORT: data32x 0 0 8 0 INPUT NODEFVAL data32x[7..0]
-- Retrieval info: USED_PORT: data33x 0 0 8 0 INPUT NODEFVAL data33x[7..0]
-- Retrieval info: USED_PORT: data34x 0 0 8 0 INPUT NODEFVAL data34x[7..0]
-- Retrieval info: USED_PORT: data35x 0 0 8 0 INPUT NODEFVAL data35x[7..0]
-- Retrieval info: USED_PORT: data36x 0 0 8 0 INPUT NODEFVAL data36x[7..0]
-- Retrieval info: USED_PORT: data37x 0 0 8 0 INPUT NODEFVAL data37x[7..0]
-- Retrieval info: USED_PORT: data38x 0 0 8 0 INPUT NODEFVAL data38x[7..0]
-- Retrieval info: USED_PORT: data39x 0 0 8 0 INPUT NODEFVAL data39x[7..0]
-- Retrieval info: USED_PORT: data3x 0 0 8 0 INPUT NODEFVAL data3x[7..0]
-- Retrieval info: USED_PORT: data40x 0 0 8 0 INPUT NODEFVAL data40x[7..0]
-- Retrieval info: USED_PORT: data41x 0 0 8 0 INPUT NODEFVAL data41x[7..0]
-- Retrieval info: USED_PORT: data42x 0 0 8 0 INPUT NODEFVAL data42x[7..0]
-- Retrieval info: USED_PORT: data43x 0 0 8 0 INPUT NODEFVAL data43x[7..0]
-- Retrieval info: USED_PORT: data44x 0 0 8 0 INPUT NODEFVAL data44x[7..0]
-- Retrieval info: USED_PORT: data45x 0 0 8 0 INPUT NODEFVAL data45x[7..0]
-- Retrieval info: USED_PORT: data46x 0 0 8 0 INPUT NODEFVAL data46x[7..0]
-- Retrieval info: USED_PORT: data47x 0 0 8 0 INPUT NODEFVAL data47x[7..0]
-- Retrieval info: USED_PORT: data48x 0 0 8 0 INPUT NODEFVAL data48x[7..0]
-- Retrieval info: USED_PORT: data49x 0 0 8 0 INPUT NODEFVAL data49x[7..0]
-- Retrieval info: USED_PORT: data4x 0 0 8 0 INPUT NODEFVAL data4x[7..0]
-- Retrieval info: USED_PORT: data50x 0 0 8 0 INPUT NODEFVAL data50x[7..0]
-- Retrieval info: USED_PORT: data51x 0 0 8 0 INPUT NODEFVAL data51x[7..0]
-- Retrieval info: USED_PORT: data52x 0 0 8 0 INPUT NODEFVAL data52x[7..0]
-- Retrieval info: USED_PORT: data53x 0 0 8 0 INPUT NODEFVAL data53x[7..0]
-- Retrieval info: USED_PORT: data54x 0 0 8 0 INPUT NODEFVAL data54x[7..0]
-- Retrieval info: USED_PORT: data55x 0 0 8 0 INPUT NODEFVAL data55x[7..0]
-- Retrieval info: USED_PORT: data56x 0 0 8 0 INPUT NODEFVAL data56x[7..0]
-- Retrieval info: USED_PORT: data57x 0 0 8 0 INPUT NODEFVAL data57x[7..0]
-- Retrieval info: USED_PORT: data58x 0 0 8 0 INPUT NODEFVAL data58x[7..0]
-- Retrieval info: USED_PORT: data59x 0 0 8 0 INPUT NODEFVAL data59x[7..0]
-- Retrieval info: USED_PORT: data5x 0 0 8 0 INPUT NODEFVAL data5x[7..0]
-- Retrieval info: USED_PORT: data60x 0 0 8 0 INPUT NODEFVAL data60x[7..0]
-- Retrieval info: USED_PORT: data61x 0 0 8 0 INPUT NODEFVAL data61x[7..0]
-- Retrieval info: USED_PORT: data62x 0 0 8 0 INPUT NODEFVAL data62x[7..0]
-- Retrieval info: USED_PORT: data63x 0 0 8 0 INPUT NODEFVAL data63x[7..0]
-- Retrieval info: USED_PORT: data64x 0 0 8 0 INPUT NODEFVAL data64x[7..0]
-- Retrieval info: USED_PORT: data65x 0 0 8 0 INPUT NODEFVAL data65x[7..0]
-- Retrieval info: USED_PORT: data66x 0 0 8 0 INPUT NODEFVAL data66x[7..0]
-- Retrieval info: USED_PORT: data67x 0 0 8 0 INPUT NODEFVAL data67x[7..0]
-- Retrieval info: USED_PORT: data68x 0 0 8 0 INPUT NODEFVAL data68x[7..0]
-- Retrieval info: USED_PORT: data69x 0 0 8 0 INPUT NODEFVAL data69x[7..0]
-- Retrieval info: USED_PORT: data6x 0 0 8 0 INPUT NODEFVAL data6x[7..0]
-- Retrieval info: USED_PORT: data70x 0 0 8 0 INPUT NODEFVAL data70x[7..0]
-- Retrieval info: USED_PORT: data71x 0 0 8 0 INPUT NODEFVAL data71x[7..0]
-- Retrieval info: USED_PORT: data72x 0 0 8 0 INPUT NODEFVAL data72x[7..0]
-- Retrieval info: USED_PORT: data73x 0 0 8 0 INPUT NODEFVAL data73x[7..0]
-- Retrieval info: USED_PORT: data74x 0 0 8 0 INPUT NODEFVAL data74x[7..0]
-- Retrieval info: USED_PORT: data75x 0 0 8 0 INPUT NODEFVAL data75x[7..0]
-- Retrieval info: USED_PORT: data76x 0 0 8 0 INPUT NODEFVAL data76x[7..0]
-- Retrieval info: USED_PORT: data77x 0 0 8 0 INPUT NODEFVAL data77x[7..0]
-- Retrieval info: USED_PORT: data78x 0 0 8 0 INPUT NODEFVAL data78x[7..0]
-- Retrieval info: USED_PORT: data79x 0 0 8 0 INPUT NODEFVAL data79x[7..0]
-- Retrieval info: USED_PORT: data7x 0 0 8 0 INPUT NODEFVAL data7x[7..0]
-- Retrieval info: USED_PORT: data80x 0 0 8 0 INPUT NODEFVAL data80x[7..0]
-- Retrieval info: USED_PORT: data81x 0 0 8 0 INPUT NODEFVAL data81x[7..0]
-- Retrieval info: USED_PORT: data82x 0 0 8 0 INPUT NODEFVAL data82x[7..0]
-- Retrieval info: USED_PORT: data83x 0 0 8 0 INPUT NODEFVAL data83x[7..0]
-- Retrieval info: USED_PORT: data84x 0 0 8 0 INPUT NODEFVAL data84x[7..0]
-- Retrieval info: USED_PORT: data85x 0 0 8 0 INPUT NODEFVAL data85x[7..0]
-- Retrieval info: USED_PORT: data86x 0 0 8 0 INPUT NODEFVAL data86x[7..0]
-- Retrieval info: USED_PORT: data87x 0 0 8 0 INPUT NODEFVAL data87x[7..0]
-- Retrieval info: USED_PORT: data88x 0 0 8 0 INPUT NODEFVAL data88x[7..0]
-- Retrieval info: USED_PORT: data89x 0 0 8 0 INPUT NODEFVAL data89x[7..0]
-- Retrieval info: USED_PORT: data8x 0 0 8 0 INPUT NODEFVAL data8x[7..0]
-- Retrieval info: USED_PORT: data90x 0 0 8 0 INPUT NODEFVAL data90x[7..0]
-- Retrieval info: USED_PORT: data91x 0 0 8 0 INPUT NODEFVAL data91x[7..0]
-- Retrieval info: USED_PORT: data92x 0 0 8 0 INPUT NODEFVAL data92x[7..0]
-- Retrieval info: USED_PORT: data93x 0 0 8 0 INPUT NODEFVAL data93x[7..0]
-- Retrieval info: USED_PORT: data94x 0 0 8 0 INPUT NODEFVAL data94x[7..0]
-- Retrieval info: USED_PORT: data95x 0 0 8 0 INPUT NODEFVAL data95x[7..0]
-- Retrieval info: USED_PORT: data96x 0 0 8 0 INPUT NODEFVAL data96x[7..0]
-- Retrieval info: USED_PORT: data97x 0 0 8 0 INPUT NODEFVAL data97x[7..0]
-- Retrieval info: USED_PORT: data98x 0 0 8 0 INPUT NODEFVAL data98x[7..0]
-- Retrieval info: USED_PORT: data99x 0 0 8 0 INPUT NODEFVAL data99x[7..0]
-- Retrieval info: USED_PORT: data9x 0 0 8 0 INPUT NODEFVAL data9x[7..0]
-- Retrieval info: USED_PORT: result 0 0 8 0 OUTPUT NODEFVAL result[7..0]
-- Retrieval info: USED_PORT: sel 0 0 8 0 INPUT NODEFVAL sel[7..0]
-- Retrieval info: CONNECT: result 0 0 8 0 @result 0 0 8 0
-- Retrieval info: CONNECT: @data 1 255 8 0 data255x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 254 8 0 data254x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 253 8 0 data253x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 252 8 0 data252x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 251 8 0 data251x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 250 8 0 data250x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 249 8 0 data249x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 248 8 0 data248x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 247 8 0 data247x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 246 8 0 data246x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 245 8 0 data245x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 244 8 0 data244x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 243 8 0 data243x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 242 8 0 data242x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 241 8 0 data241x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 240 8 0 data240x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 239 8 0 data239x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 238 8 0 data238x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 237 8 0 data237x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 236 8 0 data236x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 235 8 0 data235x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 234 8 0 data234x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 233 8 0 data233x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 232 8 0 data232x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 231 8 0 data231x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 230 8 0 data230x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 229 8 0 data229x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 228 8 0 data228x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 227 8 0 data227x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 226 8 0 data226x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 225 8 0 data225x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 224 8 0 data224x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 223 8 0 data223x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 222 8 0 data222x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 221 8 0 data221x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 220 8 0 data220x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 219 8 0 data219x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 218 8 0 data218x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 217 8 0 data217x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 216 8 0 data216x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 215 8 0 data215x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 214 8 0 data214x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 213 8 0 data213x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 212 8 0 data212x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 211 8 0 data211x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 210 8 0 data210x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 209 8 0 data209x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 208 8 0 data208x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 207 8 0 data207x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 206 8 0 data206x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 205 8 0 data205x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 204 8 0 data204x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 203 8 0 data203x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 202 8 0 data202x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 201 8 0 data201x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 200 8 0 data200x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 199 8 0 data199x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 198 8 0 data198x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 197 8 0 data197x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 196 8 0 data196x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 195 8 0 data195x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 194 8 0 data194x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 193 8 0 data193x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 192 8 0 data192x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 191 8 0 data191x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 190 8 0 data190x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 189 8 0 data189x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 188 8 0 data188x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 187 8 0 data187x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 186 8 0 data186x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 185 8 0 data185x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 184 8 0 data184x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 183 8 0 data183x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 182 8 0 data182x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 181 8 0 data181x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 180 8 0 data180x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 179 8 0 data179x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 178 8 0 data178x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 177 8 0 data177x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 176 8 0 data176x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 175 8 0 data175x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 174 8 0 data174x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 173 8 0 data173x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 172 8 0 data172x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 171 8 0 data171x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 170 8 0 data170x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 169 8 0 data169x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 168 8 0 data168x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 167 8 0 data167x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 166 8 0 data166x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 165 8 0 data165x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 164 8 0 data164x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 163 8 0 data163x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 162 8 0 data162x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 161 8 0 data161x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 160 8 0 data160x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 159 8 0 data159x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 158 8 0 data158x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 157 8 0 data157x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 156 8 0 data156x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 155 8 0 data155x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 154 8 0 data154x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 153 8 0 data153x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 152 8 0 data152x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 151 8 0 data151x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 150 8 0 data150x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 149 8 0 data149x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 148 8 0 data148x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 147 8 0 data147x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 146 8 0 data146x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 145 8 0 data145x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 144 8 0 data144x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 143 8 0 data143x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 142 8 0 data142x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 141 8 0 data141x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 140 8 0 data140x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 139 8 0 data139x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 138 8 0 data138x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 137 8 0 data137x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 136 8 0 data136x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 135 8 0 data135x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 134 8 0 data134x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 133 8 0 data133x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 132 8 0 data132x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 131 8 0 data131x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 130 8 0 data130x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 129 8 0 data129x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 128 8 0 data128x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 127 8 0 data127x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 126 8 0 data126x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 125 8 0 data125x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 124 8 0 data124x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 123 8 0 data123x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 122 8 0 data122x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 121 8 0 data121x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 120 8 0 data120x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 119 8 0 data119x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 118 8 0 data118x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 117 8 0 data117x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 116 8 0 data116x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 115 8 0 data115x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 114 8 0 data114x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 113 8 0 data113x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 112 8 0 data112x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 111 8 0 data111x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 110 8 0 data110x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 109 8 0 data109x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 108 8 0 data108x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 107 8 0 data107x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 106 8 0 data106x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 105 8 0 data105x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 104 8 0 data104x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 103 8 0 data103x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 102 8 0 data102x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 101 8 0 data101x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 100 8 0 data100x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 99 8 0 data99x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 98 8 0 data98x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 97 8 0 data97x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 96 8 0 data96x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 95 8 0 data95x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 94 8 0 data94x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 93 8 0 data93x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 92 8 0 data92x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 91 8 0 data91x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 90 8 0 data90x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 89 8 0 data89x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 88 8 0 data88x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 87 8 0 data87x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 86 8 0 data86x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 85 8 0 data85x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 84 8 0 data84x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 83 8 0 data83x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 82 8 0 data82x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 81 8 0 data81x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 80 8 0 data80x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 79 8 0 data79x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 78 8 0 data78x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 77 8 0 data77x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 76 8 0 data76x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 75 8 0 data75x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 74 8 0 data74x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 73 8 0 data73x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 72 8 0 data72x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 71 8 0 data71x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 70 8 0 data70x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 69 8 0 data69x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 68 8 0 data68x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 67 8 0 data67x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 66 8 0 data66x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 65 8 0 data65x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 64 8 0 data64x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 63 8 0 data63x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 62 8 0 data62x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 61 8 0 data61x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 60 8 0 data60x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 59 8 0 data59x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 58 8 0 data58x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 57 8 0 data57x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 56 8 0 data56x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 55 8 0 data55x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 54 8 0 data54x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 53 8 0 data53x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 52 8 0 data52x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 51 8 0 data51x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 50 8 0 data50x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 49 8 0 data49x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 48 8 0 data48x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 47 8 0 data47x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 46 8 0 data46x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 45 8 0 data45x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 44 8 0 data44x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 43 8 0 data43x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 42 8 0 data42x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 41 8 0 data41x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 40 8 0 data40x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 39 8 0 data39x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 38 8 0 data38x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 37 8 0 data37x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 36 8 0 data36x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 35 8 0 data35x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 34 8 0 data34x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 33 8 0 data33x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 32 8 0 data32x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 31 8 0 data31x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 30 8 0 data30x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 29 8 0 data29x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 28 8 0 data28x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 27 8 0 data27x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 26 8 0 data26x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 25 8 0 data25x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 24 8 0 data24x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 23 8 0 data23x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 22 8 0 data22x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 21 8 0 data21x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 20 8 0 data20x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 19 8 0 data19x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 18 8 0 data18x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 17 8 0 data17x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 16 8 0 data16x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 15 8 0 data15x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 14 8 0 data14x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 13 8 0 data13x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 12 8 0 data12x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 11 8 0 data11x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 10 8 0 data10x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 9 8 0 data9x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 8 8 0 data8x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 7 8 0 data7x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 6 8 0 data6x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 5 8 0 data5x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 4 8 0 data4x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 3 8 0 data3x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 2 8 0 data2x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 1 8 0 data1x 0 0 8 0
-- Retrieval info: CONNECT: @data 1 0 8 0 data0x 0 0 8 0
-- Retrieval info: CONNECT: @sel 0 0 8 0 sel 0 0 8 0
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX_REG.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX_REG.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX_REG.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX_REG.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MUX_REG_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
